.subckt MLP ACTIVATIONPREV TARGET ACTIVATIONNEXT1 ACTIVATIONNEXT2 XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUTTARGET1L OUTPUTTARGET1R OUTPUTTARGET2L OUTPUTTARGET2R

#need Oi.T + Oi.!Oj + T.!Oj
#delays so timing matches up
Xactdelayed DELAY7 ACTIVATIONPREV  XIN1 B6 XIN2 A5 DCIN DC6  0 DELAYOUTACT1  0 DELAYOUTACT2
XTARGETdelayed DELAY7 TARGET  B6 B7 A5 A6 DC6 DC7 0 DELAYOUTTARGET1  0 DELAYOUTTARGET2 

#Oi.T - correct
Xand1  AND A6 A7 B7 B8 DELAYOUTTARGET1 DELAYOUTACT1 DC7 DC8 andout1
#Oi.Oj! - correct
Xand2  AND A7 A8 B8 B9 DELAYOUTACT2 ACTIVATIONNEXT1 DC8 DC9 andout2
#T.Oj - correct
Xand3  AND A8 A9 B9 B10 DELAYOUTTARGET2 ACTIVATIONNEXT2 DC9 DC10 andout3

#MLP : D = Oi.T + Oi.!Oj + T.!Oj - correct
X3OR OR3 XOUT2 A9 XOUT1 B10  ANDOUT1 ANDOUT2 ANDOUT3 DC10 DCOUT OUTPUTTARGET1L OUTPUTTARGET1R OUTPUTTARGET2L OUTPUTTARGET2R

.ends MLP



#3-input AND gate

.subckt AND3 XIN1 XOUT1 XIN2 XOUT2 DINA DINB DIND DCIN DCOUT DOUT1 DOUT2

#AND so C=0
vINC INconst1 0 PWL(0 0 1ps -5mV 200ps -5mV 400ps -5mV 401ps -5mV 600ps -5mV )
RIN3    INconst1   INconst2   1000
LIN3    INconst2   DINC   0.1p
***********buffer1********

#INDUCTANCES
K1_1 L1_X L1_D 0.2322
K1_2 L1_D L1_OUT 3.27E-5
K1_3 L1_X L1_OUT 3.68E-5
K1_4 L1_D L1_Q 4.9E-4
K1_5 L1_X L1_Q 5.11E-4
K1_6 L1_OUT L1_Q -0.15
K1_7 L1_2 L1_D -0.1556
K1_8 L1_2 L1_X -0.228
K1_9 L1_X L1_1 -0.2284
K1_10 L1_D L1_1 -0.1559


L1_1 A_LEFT A 1.51p
L1_2 A A_RIGHT 1.51p
L1_D DCIN DC4 6.94p
#was 6.94p
L1_IN DINA A 1.526p
L1_OUT 0 BUFFIN  25.3p
L1_Q A 0 5.84p
#was 5.84
L1_X XIN1 XLINE1 6.51p

B1_1 A_LEFT 0 11 jjmit area=0.5
B1_2 A_RIGHT 0 12 jjmit area=0.5

***********buffer2********

K2_1 L2_X L2_D 0.2322
K2_2 L2_D L2_OUT 3.27E-5
K2_3 L2_X L2_OUT 3.68E-5
K2_4 L2_D L2_Q 4.9E-4
K2_5 L2_X L2_Q 5.11E-4
K2_6 L2_OUT L2_Q -0.15
K2_7 L2_2 L2_D -0.1556
K2_8 L2_2 L2_X -0.228
K2_9 L2_X L2_1 -0.2284
K2_10 L2_D L2_1 -0.1559


L2_1 B_LEFT B 1.51p
L2_2 B B_RIGHT 1.51p
L2_D DC4 DC5 6.94p
#was 6.94p
L2_IN DINB B 1.526p
L2_OUT  0 BUFFIN  25.3p
L2_Q B 0 5.84p
#was 5.84
L2_X XLINE1 XLINE2 6.51p

B2_1 B_LEFT 0 13 jjmit area=0.5
B2_2 B_RIGHT 0 14 jjmit area=0.5

***********buffer3********

K3_1 L3_X L3_D 0.2322
K3_2 L3_D L3_OUT 3.27E-5
K3_3 L3_X L3_OUT 3.68E-5
K3_4 L3_D L3_Q 4.9E-4
K3_5 L3_X L3_Q 5.11E-4
K3_6 L3_OUT L3_Q -0.3878
K3_7 L3_2 L3_D -0.1556
K3_8 L3_2 L3_X -0.228
K3_9 L3_X L3_1 -0.2284
K3_10 L3_D L3_1 -0.1559


L3_1 C_LEFT C 1.51p
L3_2 C C_RIGHT 1.51p
L3_D DC5 DC6 6.94p
#was 6.94p
L3_IN DINC C 1.526p
L3_OUT  0 BUFFIN  25.3p
L3_Q C 0 5.84p
#was 5.84
L3_X XLINE2 XLINE3 6.51p

B3_1 C_LEFT 0 15 jjmit area=0.5
B3_2 C_RIGHT 0 16 jjmit area=0.5

***********buffer4********

K4_1 L4_X L4_D 0.2322
K4_2 L4_D L4_OUT 3.27E-5
K4_3 L4_X L4_OUT 3.68E-5
K4_4 L4_D L4_Q 4.9E-4
K4_5 L4_X L4_Q 5.11E-4
K4_6 L4_OUT L4_Q -0.15
K4_7 L4_2 L4_D -0.1556
K4_8 L4_2 L4_X -0.228
K4_9 L4_X L4_1 -0.2284
K4_10 L4_D L4_1 -0.1559


L4_1 D_LEFT D 1.51p
L4_2 D D_RIGHT 1.51p
L4_D DC6 DC7 6.94p
#was 6.94p
L4_IN DIND D 1.526p
L4_OUT  0 BUFFIN  25.3p
L4_Q D 0 5.84p
#was 5.84
L4_X XLINE3 XOUT1 6.51p

B4_1 D_LEFT 0 15D jjmit area=0.5
B4_2 D_RIGHT 0 16D jjmit area=0.5



***********buffer OUT ********

K5_1 L5_X L5_D 0.2322
K5_2 L5_D L5_OUT1 3.27E-5
K5_3 L5_X L5_OUT1 3.68E-5
K5_4 L5_D L5_Q 4.9E-4
K5_5 L5_X L5_Q 5.11E-4
K5_6 L5_OUT1 L5_Q -0.3878
K5_7 L5_2 L5_D -0.1556
K5_8 L5_2 L5_X -0.228
K5_9 L5_X L5_1 -0.2284
K5_10 L5_D L5_1 -0.1559
K5_11 L5_OUT2 L5_Q -0.3878
K5_12 L5_D L5_OUT2 3.27E-5
K5_13 L5_X L5_OUT2 3.68E-5

#tinkered with l4q which was 0.14p now 1.514 may change back to 5.14p
L5_1 OUT_LEFT OUT 1.51p
L5_2 OUT OUT_RIGHT 1.51p
L5_D DCOUT DC7 6.94p
#was 6.94p
L5_IN BUFFIN OUT 1.526p
L5_OUT1  0 DOUT1  25.3p
L5_OUT2  0 DOUT2  25.3p
L5_Q OUT 0 8.84p
#was 13.84
#ADJUST TO CHANGE OUTPUT WAVEFORM
L5_X XIN2 XOUT2 6.51p

B5_1 OUT_LEFT 0 17 jjmit area=0.5
B5_2 OUT_RIGHT 0 18 jjmit area=0.5
.ends and3
#CKT TO TRASMIT PULSE TO NEXT SYNAPSE
.subckt TRANSMIT INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT DCCIN DCCOUT OUTPUT

XBUFF bfrconv XIN1 INPUT XOUT1 DCOUT DCIN DOUTLBUFF 0
XCONV AQFP2RSFQ3 XOUT2 XIN2 DOUTLBUFF RSFQOUT  DCCIN DCCOUT

#TRANSMISISON STAGE
#SPLITTING
XSPLIT MULTISPLIT RSFQOUT SPLIT1 SPLIT2 SPLIT3 SPLIT4 SPLIT5 SPLIT6 SPLIT7 SPLIT8
#CURRENT PULSES
#FIRST ACTIVATION
XDC1 DCPULSER SPLIT1 DCOUT1
XDC2 DCPULSER SPLIT2 DCOUT2
XDC3 DCPULSER SPLIT3 DCOUT3 
XDC4 DCPULSER SPLIT4 DCOUT4 
XDC5 DCPULSER SPLIT5 DCOUT5 
XDC6 DCPULSER SPLIT6 DCOUT6 
XDC7 DCPULSER SPLIT7 DCOUT7
XDC8 DCPULSER SPLIT8 DCOUT8
.PARAM ROUT=0.7
rOUT1 DCOUT1 OUTPUT ROUT
rOUT2 DCOUT2 OUTPUT ROUT
rOUT3 DCOUT3 OUTPUT ROUT
rOUT4 DCOUT4 OUTPUT ROUT
rOUT5 DCOUT5 OUTPUT ROUT
rOUT6 DCOUT6 OUTPUT ROUT
rOUT7 DCOUT7 OUTPUT ROUT
rOUT8 DCOUT8 OUTPUT ROUT

.ends TRANSMIT
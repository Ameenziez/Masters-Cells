.subckt COMP4 XIN DIN XOUT DCIN DCOUT DOUTL1 DOUTR1 DOUTL2 DOUTR2 DOUTL3 DOUTR3 DOUTL4 DOUTR4  CONST
B1 8 0 11 jjmit area=0.5
B2 9 0 12 jjmit area=0.5
K1 LX LD 0.2322
K2 LD LOUT1 3.27E-5
K3 LX LOUT1 3.68E-5
K4 LD LQ 4.9E-4
K5 LX LQ 5.11E-4
K6 LOUT1 LQ -0.28
K7 L2 LD -0.1556
K8 L2 LX -0.228
K9 LX L1 -0.2284
K10 LD L1 -0.15559
K11 LD LOUT2 3.27E-5
K12 LX LOUT2 3.68E-5
K13 LOUT2 LQ -0.28
K14 LD LOUT3 3.27E-5
K15 LX LOUT3 3.68E-5
K16 LOUT3 LQ -0.28
K17 LD LOUT4 3.27E-5
K18 LX LOUT4 3.68E-5
K19 LOUT4 LQ -0.28


#iconst 0 CONST PWL(0 0 20p 45u)
#CHANGEWD COMP CIRCUIT TO HAVE CONST INPUT TO SUBCKT (11'S VERSION DIDNT HAVE THI ALREADY...)
#45 WORKS CURRENT CONFIG
Lconst CONST 0 20p
Lconstout 7Q 7 25.5P
Kconst  Lconst Lconstout 0.1
L1 8 7 1.51p
L2 7 9 1.51p
LD DCIN DCOUT 7.94p
#was 7.94p
LIN DIN 7Q 1.526p
LOUT1 DOUTL1 DOUTR1 25.3p

LOUT2 DOUTL2 DOUTR2 25.3p
LOUT3 DOUTL3 DOUTR3 25.3p
LOUT4 DOUTL4 DOUTR4 25.3p
LQ 7 0 5.84p
#WAS 5.84
LX XIN XOUT 6.51p
.ends COMP4

.subckt COMP4F XIN DIN XOUT DCIN DCOUT DOUTL1 DOUTR1 DOUTL2 DOUTR2 DOUTL3 DOUTR3 DOUTL4 DOUTR4 CONST
B1 8 0 11 jjmit area=0.5
B2 9 0 12 jjmit area=0.5
K1 LX LD 0.2322
K2 LD LOUT1 3.27E-5
K3 LX LOUT1 3.68E-5
K4 LD LQ 4.9E-4
K5 LX LQ 5.11E-4
K6 LOUT1 LQ -0.28
K7 L2 LD -0.1556
K8 L2 LX -0.228
K9 LX L1 -0.2284
K10 LD L1 -0.15559
K11 LD LOUT2 3.27E-5
K12 LX LOUT2 3.68E-5
K13 LOUT2 LQ -0.28
K14 LD LOUT3 3.27E-5
K15 LX LOUT3 3.68E-5
K16 LOUT3 LQ -0.28
K17 LD LOUT4 3.27E-5
K18 LX LOUT4 3.68E-5
K19 LOUT4 LQ -0.28
K20 LD LOUT5 3.27E-5
K21 LX LOUT5 3.68E-5
K22 LOUT5 LQ -0.2


#iconst 0 CONST PWL(0 0 20p 45u)
#CHANGEWD COMP CIRCUIT TO HAVE CONST INPUT TO SUBCKT (11'S VERSION DIDNT HAVE THI ALREADY...)
#45 WORKS CURRENT CONFIG
Lconst CONST 0 20p
Lconstout 7Q 7 25.5P
Kconst  Lconst Lconstout 0.1
L1 8 7 1.51p
L2 7 9 1.51p
LD DCIN DCOUT 7.94p
#was 7.94p
LIN DIN 7Q 1.526p
LOUT1 DOUTL1 DOUTR1 25.3p

LOUT2 DOUTL2 DOUTR2 25.3p
LOUT3 DOUTL3 DOUTR3 25.3p
LOUT4 DOUTL4 DOUTR4 25.3p
LOUT5 DOUTL5 DOUTR5 25.3p
LQ 7 0 5.84p
#WAS 5.84
LX XIN XOUT 6.51p
RSHUNT 8 0 100
.ends COMP4F


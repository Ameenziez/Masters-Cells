

.subckt PERCEPTRON2LAYER XIN1 XOUT1 XIN2 XOUT2 INPUT ACTIVATIONP ACTIVATIONN TARGET DCIN DCOUT INCR DECR

XINPUT bfrsplit2 XIN1 INPUT X1LINE1 DCIN DC5  DOUTRIN 0 DOUTRIN2 0
XTARGET bfrsplit4 X1LINE1 TARGET X1LINE2 DC5 DC6 DOUTRT1 0 0 DOUTLT2 DOUTLT3 0 DOUTLT4 0

XDECR AND3R     X2LINE1  XIN2 X1LINE2 X1LINE3 DOUTRIN ACTIVATIONN DOUTRT1   DC7 DC6  DECR 0
XINCR AND3R     XOUT2  X2LINE1 X1LINE3 XOUT1 DOUTRIN2 ACTIVATIONP DOUTLT2   DCOUT DC7  INCR 0

#XINPUT0 bfr XIN1 INPUT X1LINE1 DCIN DC5 DOUTIN 0
#XINPUT bfrsplit2 XIN2 DOUTIN X2LINE1 DC6 DC5  DOUTRIN 0 DOUTRIN2 0
#XTARGET0 bfr X1LINE1 TARGET X1LINE2 DC6 DC7 0 TARGETIN 
#XTARGET bfrsplit4 X2LINE1 TARGETIN X2LINE2 DC8 DC7 DOUTRT1 0 0 DOUTLT2 DOUTLT3 0 DOUTLT4 0


#XDECR AND3R     X1LINE3 X1LINE2  X2LINE3  X2LINE2  DOUTRIN ACTIVATIONN DOUTRT1   DC9 DC8   DECR 0
#XINCR AND3R     XOUT1  X1LINE3 XOUT2 X2LINE3  DOUTRIN2 ACTIVATIONP DOUTLT2   DCOUT DC9 INCR 0

#FLIPPED ALL CLKS AND DC

.ends PERCEPTRON2LAYER




.subckt PERCEPTRON2LAYER2 XIN1 XOUT1 XIN2 XOUT2 INPUT ACTIVATIONP ACTIVATIONN TARGET DCIN DCOUT INCR DECR

XINPUT bfrsplit2 XIN1 INPUT X1LINE1 DCIN DC5  DOUTRIN 0 DOUTRIN2 0
XTARGET bfrsplit2 X1LINE1 TARGET X1LINE2 DC5 DC6 DOUTRT1 0 0 DOUTLT2 

XDECR AND3R     X2LINE1  XIN2 X1LINE2 X1LINE3 DOUTRIN ACTIVATIONN DOUTRT1   DC7 DC6  DECR 0
XINCR AND3R     XOUT2  X2LINE1 X1LINE3 XOUT1 DOUTRIN2 ACTIVATIONP DOUTLT2   DCOUT DC7  INCR 0

#XINPUT0 bfr XIN1 INPUT X1LINE1 DCIN DC5 DOUTIN 0
#XINPUT bfrsplit2 XIN2 DOUTIN X2LINE1 DC6 DC5  DOUTRIN 0 DOUTRIN2 0
#XTARGET0 bfr X1LINE1 TARGET X1LINE2 DC6 DC7 0 TARGETIN 
#XTARGET bfrsplit4 X2LINE1 TARGETIN X2LINE2 DC8 DC7 DOUTRT1 0 0 DOUTLT2 DOUTLT3 0 DOUTLT4 0


#XDECR AND3R     X1LINE3 X1LINE2  X2LINE3  X2LINE2  DOUTRIN ACTIVATIONN DOUTRT1   DC9 DC8   DECR 0
#XINCR AND3R     XOUT1  X1LINE3 XOUT2 X2LINE3  DOUTRIN2 ACTIVATIONP DOUTLT2   DCOUT DC9 INCR 0

#FLIPPED ALL CLKS AND DC

.ends PERCEPTRON2LAYER2

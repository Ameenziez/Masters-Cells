.SUBCKT CONV CLKIN CLKOUT DCIN DCOUT AQFPP AQFPM INCR DECR
XCONVP AQFP2RSFQ A6 CLKIN AQFPP RSFQOUTP DC6 DCIN
XCONVM AQFP2RSFQ CLKOUT A6 AQFPM RSFQOUTM DCOUT DC6
#was 5ohms,1p - works with 5, 30p for some reason
#TTESTP    RSFQOUTP         0          RSFQOUTPT          0  Z0=5 TD=30p
#TTESTM    RSFQOUTM         0          RSFQOUTMT          0  Z0=5 TD=30p
RCONN1 RSFQOUTP RSFQOUTPT 1
RCONN2 RSFQOUTM RSFQOUTMT 1 
XBUFF1 LSmitll_bufft  RSFQOUTPT INCR
XBUFF2 LSmitll_bufft  RSFQOUTMT DECR
.ends CONV

#works well!
#got the data to propagate
.include LSmitll_DCSFQ_PTLTX_v1p5.cir
.include LSmitll_bufft_v1p5.cir
.include LSmitll_PTLRX_SFQDC_v1p5.cir
.include LSmitll_SPLITT_v1p5.cir
.INCLUDE LSMITLL_JTLT_V1P5.CIR
.INCLUDE LSMITLL_MERGET_V1P5.CIR
.include storeedit.cir
.INCLUDE COMPONENTSEDIT.CIR
.INCLUDE COMP3.CIR
.INCLUDE COMP4.CIR
.INCLUDE COMP5.CIR
.INCLUDE COMP6.CIR
.include conv.cir
.INCLUDE synapsenext2.CIR
.INCLUDE DCPULSER.CIR
.INCLUDE MULTISPLIT.CIR
.include transmit.cir
.INCLUDE DELAY7.CIR
.INCLUDE AND.CIR
.INCLUDE AND3.CIR
.INCLUDE OR3.CIR
.include PERCEPTRON.CIR
.include PERCEPTRON2.CIR
.include CONVINTERFACE.cir


# TRY SHIFTING CLK OF OUTPUT BACK A BIT...

.tran 1ps 25000PS 0ps 1p
#MLP:
#D=Oi.T + Oi.!Oj + T.!Oj 

#setup circuitry
VAC1   A1   0   SIN(0 723mV 10GHz 200Ps 0)
RAC1   A1   A2   1000
LAC1   A2   A3   0.1p
VAC2   B1   0   SIN(0 723mV 10GHz 175.0ps 0)
RAC2   B1   B2   1000
LAC2   B2   B3   0.1p
VDC    DC1   0   pwl(0 0 20p 1023mV)
RDC    DC1   DC2   1000
LDC    DC2   DC3  0.1p
VDCconv    DCc1   0   PWL(0ps 0mV 20ps 1023mV 1.881e-08 1023mV 1.8811000000000002e-08 0)
RDCconv    DCc1   DCc2  640
LDCconv    DCc2   DCc3   0.1p




#SECOND LAYER SYNAPSE 1
IINITAL21 0 INITIAL21 PWL( 0 0 20P flx21*2*22.6U)
XSTORE21 BISTORE SFQOUTPLUS21 SFQOUTMINUS21 WEIGHTL21 WEIGHTR21


#NEXT LAYER BIAS
#Iactualsynbias21 0 ACTUALSYNB21x PWL(0 0 640P 0 665P 670U 700P 0 840P 0 865P 670U 900P 0  1040P 0 1065P 670U 1100P 0 1240P 0 1265P 670U 1300P 0  )
LSYNB21 ACTUALSYNB21x ACTUALSYNB21 1p  
KSYNB21 LSYNB21 LSYNADJUSTB21 0.3
LSYNADJUSTB21 0 ADJUSTB21 5P 

#SPLIT TARGET BETWEEN 2 NEURONS
LTARGET1 TARGET0 TARGET1 1p
LTARGET2 TARGET0 TARGET2 1p

#SPLIT INPUTS BETWEEN 2 NEURONS
LINPUT1 IN1 INPUT11 1P
LINPUT2 IN1 INPUT12 1P
LINPUT3 IN2 INPUT13 1P
LINPUT4 IN2 INPUT14 1P
LINPUTBIAS11 INB11 INPUTB12 1P
LINPUTBIAS12 INB11 INPUTB13 1P


IINITALB21 0 INITIALB21 PWL( 0 0 20P flxb21*2*22.6U)
XSTOREB21 BISTORE SFQOUTPLUSB21 SFQOUTMINUSB21 WEIGHTLB21 WEIGHTRB21

X21 SYNAPSEfastestnext2 OUTPUTAXON DOUT22 DOUT21  WEIGHTL21 WEIGHTR21 INITIAL21
XB21 SYNAPSEfastestnext2 ACTUALSYNB21  0 DOUT23   WEIGHTLB21 WEIGHTRB21 INITIALB21

.param flx11 = -2
.param flx12 = 2
.param flx13 = 3
.param flx14 = 0
.param flxb11 = 1
.param flxb12 = -1
.param flx21 = -4
.param flx22 = 3
.param flxb21 = 0


IINITAL11 0 INITIAL11 PWL( 0 0 20P -22U*2*flx11)
IINITAL12 0 INITIAL12 PWL( 0 0 20P -22u*2*flx12)
IINITALB11 0 INITIALB11 PWL( 0 0 20P -22u*2*flxb11)

IINITAL13 0 INITIAL13 PWL( 0 0 20P -22U*2*flx13)
IINITAL14 0 INITIAL14 PWL( 0 0 20P -22u*2*flx14)
IINITALB12 0 INITIALB12 PWL( 0 0 20P -22u*flxb12)


##FINAL ACTIVATION - this works 
#ITHRESH11 0 THRESH11 PWL(0 0 20p 200U)
#ITHRESH12 0 THRESH12 PWL(0 0 20p 18U)
#ITHRESH21 0 THRESH21 PWL(0 0 20p -20U)
ITHRESH11 0 THRESH11 PWL(0 0 20p 195U)
ITHRESH12 0 THRESH12 PWL(0 0 20p 175U)
ITHRESH21 0 THRESH21 PWL(0 0 20p -5U)
#was like 23u
XACTfinal COMP6 A5 DOUT21 A6  DC6 DC5   DOUTFINAL1 0   DOUTFINAL2 0   DOUTFINAL3 0   DOUTFINAL4  0 DOUTFINAL5 0 DOUTFINAL6 0   THRESH21

XNEURON1 3NEURON2 INPUT11 INPUT13 INPUTB12 TARGET1 DOUTFINAL1 DOUTFINAL2 THRESH11 A3 A5 B3 B4 DC3 DC5 DCC3 DCC4  OUTPUT1 0    OUTPUT2 0 OUTPUTAXON 0 DELAYEDTARGETP  0 DELAYEDTARGETN 0 DELAYEDTARGETP2   INITIAL11 INITIAL12 INITIALB11
          #x3NEURON2 INPUT1 INPUT2 INPUTBIAS TARGET DOUTFINAL1 DOUTFINAL2 THRESH XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT DCCIN DCCOUT OUTPUT OUTPUTAXON

xbfrout1 bfrsplit4 B4 DOUTFINAL3 B6 dc6 DC8  0 actfinaloutp actfinaloutn 0 0 actfinaloutp2  actfinaloutn2 0 


#XPERCEPTRON21 PERCEPTRON   B6  B7 A7 A6   OUTPUT1  actfinaloutp actfinaloutn DELAYEDTARGETP   DC8 DC9 INCR21 DECR21
XPERCEPTRON21 PERCEPTRON2LAYER   B6  B7 A7 A6   OUTPUT1  actfinaloutp actfinaloutn DELAYEDTARGETP   DC8 DC9 INCR21 DECR21
XCONVO CONV A7 A8   DCC5 DCC4  INCR21 DECR21 SFQOUTPLUS21 SFQOUTMINUS21

#XPERCEPTRONb21 PERCEPTRON   B7  B8 A9 A8   ADJUSTB21  actfinaloutp2 actfinaloutn2 DELAYEDTARGETP2   DC9 DC10 INCRb21 DECRb21
XPERCEPTRONb21 PERCEPTRON2LAYER   B7  B8 A9 A8   ADJUSTB21  actfinaloutp2 actfinaloutn2 DELAYEDTARGETP2   DC9 DC10 INCRb21 DECRb21

XCONVb21 CONV A9 A10   DCC6 DCC5  INCRb21 DECRb21 SFQOUTPLUSb21 SFQOUTMINUSb21

XNEURON2 3NEURON2 INPUT12 INPUT14 INPUTB13 TARGET2 DOUTFINAL5 DOUTFINAL6 THRESH12 A10 A11 B8 B9 DC10 DC11 DCC6 DCC7 OUTPUT3 0  OUTPUT4 0 OUTPUTAXON2 0 DELAYEDTARGETP12  0 DELAYEDTARGETN12  DELAYEDTARGETP13  0 INITIAL13 INITIAL14 INITIALB12
IINITAL22 0 INITIAL22 PWL( 0 0 20P flx22*2*22.6U)
XSTORE22 BISTORE SFQOUTPLUS22 SFQOUTMINUS22 WEIGHTL22 WEIGHTR22


X22 SYNAPSEfastestnext2 OUTPUTAXON2 DOUT23 DOUT22  WEIGHTL22 WEIGHTR22 INITIAL22
xbfrout2 bfrsplit2 B9 DOUTFINAL4 B10 DC11 DC12  actfinaloutp3 0 0 actfinaloutn3 
#XPERCEPTRON22 PERCEPTRON   B10  0 A12 A11   OUTPUT3  actfinaloutp3 actfinaloutn3 DELAYEDTARGETP12   DC12 0 INCR22 DECR22
XPERCEPTRON22 PERCEPTRON2LAYER   B10  0 A12 A11   OUTPUT3  actfinaloutp3 actfinaloutn3 DELAYEDTARGETP2   DC12 0 INCR22 DECR22

XCONVO22 CONV A12 0   0 DCC7  INCR22 DECR22 SFQOUTPLUS22 SFQOUTMINUS22







.PRINT DEVII IIN1
.PRINT DEVII IIN2
#.print devii IINBIAS1
.PRINT DEVII ITARGET
#.print devii Iactualsynbias21
#.print devii Iactualsynbias21
#.print phase lstore1.x11.XNEURON1
#.print phase lstore1.x12.XNEURON1
#.print phase lstore1.xb11.XNEURON1
#.print phase lstore1.xb11.XNEURON2
#.print phase lq.x11.xNEURON1
#.print phase lq.x12.xNEURON1
.PRINT PHASE LQ.XACT11.XNEURON1
.PRINT PHASE LQ.XACT11.XNEURON2


#.PRINT PHASE LQ.X21
#.print phase lstore1.X21
.PRINT PHASE LSTORE1.X22
#.print phase lstore1.Xb21


#.print phase lq.XTARGET.XPERCEPTRONb21
#.print phase L1_Q.xINCR.XPERCEPTRONb21
#.print phase L2_Q.xINCR.XPERCEPTRONb21
#.print phase L4_Q.xINCR.XPERCEPTRONb21
#.print phase L5_Q.xINCR.XPERCEPTRONb21
#.print phase L1_Q.xDECR.XPERCEPTRON21
#.print phase L2_Q.xDECR.XPERCEPTRON21
#.print phase L4_Q.xDECR.XPERCEPTRON21
#.print phase L5_Q.xDECR.XPERCEPTRON21
#.print phase L1_Q.xDECR.XPERCEPTRON22
#.print phase L2_Q.xDECR.XPERCEPTRON22
#.print phase L4_Q.xDECR.XPERCEPTRON22
#.print phase L5_Q.xDECR.XPERCEPTRON22

#.print phase lq.XB21

#.print phase lq.XINPUT.XPERCEPTRONb11.xNEURON1
#.print phase lq.XTARGET.XPERCEPTRONb11.xNEURON1
#.print phase L1_Q.xINCR.XPERCEPTRONB11.xNEURON1
#.print phase L2_Q.xINCR.XPERCEPTRONB11.xNEURON1
#.print phase L4_Q.xINCR.XPERCEPTRONb11.xNEURON1
#.print phase L5_Q.xINCR.XPERCEPTRONb11.xNEURON1

#.print phase lq.XINPUT.XPERCEPTRONb11.xNEURON1
#.print phase lq.XTARGET.XPERCEPTRONb11.xNEURON1
#.print phase L1_Q.xdeCR.XPERCEPTRONB11.xNEURON1
#.print phase L2_Q.xdeCR.XPERCEPTRONB11.xNEURON1
#.print phase L4_Q.xdeCR.XPERCEPTRONb11.xNEURON1
#.print phase L5_Q.xdeCR.XPERCEPTRONb11.xNEURON1

#.print devii Iactualsynbias21
.print phase lq.XINPUT.XPERCEPTRON22
.print phase lq.XTARGET.XPERCEPTRON21
.print phase lq.XTARGET.XPERCEPTRON22
.print phase L1_Q.xINCR.XPERCEPTRON22
.print phase L2_Q.xINCR.XPERCEPTRON22
.print phase L4_Q.xINCR.XPERCEPTRON22
.print phase L5_Q.xINCR.XPERCEPTRON22
.print phase L1_Q.xdeCR.XPERCEPTRON22
.print phase L2_Q.xdeCR.XPERCEPTRON22
.print phase L4_Q.xdeCR.XPERCEPTRON22
.print phase L5_Q.xdeCR.XPERCEPTRON22
#.print phase L2_Q.xINCR.XPERCEPTRON21
#.print phase L2_Q.xINCR.XPERCEPTRONb21
#.print phase L5_Q.xINCR.XPERCEPTRON22
#.print phase L1_Q.xDECR.XPERCEPTRONb21
#.print phase L2_Q.xDECR.XPERCEPTRONb21
.print phase L4_Q.xDECR.XPERCEPTRONb21
#.print phase L5_Q.xDECR.XPERCEPTRONb21



#.PRINT DEVII ITARGET
.PRINT PHASE LQ.XACTfinal
#.PRINT PHASE LQ.XACT11.XNEURON1
#.print phase L1_Q.X3OR.XMLP.XNEURON1
#.print phase L2_Q.X3OR.XMLP.XNEURON1
#.print phase L4_Q.X3OR.XMLP.XNEURON1
#.print nodep OUTPUTTARGET3L.XNEURON1
#.print nodep OUTPUTTARGET2L.XNEURON1
#.print nodep OUTPUTTARGET1L.XNEURON1

.print phase LQ.XDELAY15.XDELAYTARGET2.XNEURON1

.SUBCKT 3NEURON2 INPUT1 INPUT2 INPUTBIAS TARGET ACTNEXT1 ACTNEXT2 THRESH XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT DCCIN DCCOUT OUTPUT1 OUTPUT1GND OUTPUT2 OUTPUT2GND OUTPUTAXON DELAYOUTTARGET3 DELAYOUTTARGET3GND DELAYOUTTARGET4 DELAYOUTTARGET4GND DELAYOUTTARGET5 DELAYOUTTARGET5GND INITIAL11 INITIAL12 INITIALB11

#INPUTS
LSYN11 INPUT1 SYN11 1p  
LSYN12 INPUT2 SYN12 1p  
LSYNB11 INPUTBIAS SYNB11 1p  
LTARGET1 TARGET TARGET1 1p
LTARGET2 TARGET1 0 1p

#COUPLINGS
KSYN11 LSYN11 LSYNADJUST11 -0.05
KSYN12 LSYN12 LSYNADJUST12 -0.05
KSYNB11 LSYNB11 LSYNADJUSTB11 -0.05
KT1 LTARGET1 LADJUSTTARGET1 -0.05
KT2 LTARGET2 LADJUSTTARGET2 -0.05
LSYNADJUST11 0 ADJUST11 5P 
LSYNADJUST12 0 ADJUST12 5P 
LSYNADJUSTB11 0 ADJUSTB11 5P 
LADJUSTTARGET1 0 ADJUSTTARGET1 5P
LADJUSTTARGET2 0 ADJUSTTARGET2 5P


#SYNAPSE 1
#IINITAL11 0 INITIAL11 PWL( 0 0 20P -80U)
XSTORE11 BISTORE SFQOUTPLUS11 SFQOUTMINUS11 WEIGHTL11 WEIGHTR11
X11 SYNAPSEfastest SYN11 DOUT12 DOUT11 WEIGHTL11 WEIGHTR11 INITIAL11
#l111 SFQOUTPLUS11 0 1p
#l112 SFQOUTMINUS11 0 1p

#SYNAPSE 2
#IINITAL12 0 INITIAL12 PWL( 0 0 20P -80U)
XSTORE12 BISTORE SFQOUTPLUS12 SFQOUTMINUS12 WEIGHTL12 WEIGHTR12
X12 SYNAPSEfastest SYN12 DOUT13 DOUT12 WEIGHTL12 WEIGHTR12 INITIAL12
#l121 SFQOUTPLUS12 0 1p
#l122 SFQOUTMINUSB12 0 1p

#SYNAPSE BIAS
#IINITALB11 0 INITIALB11 PWL( 0 0 20P -80U)
XSTOREB11 BISTORE SFQOUTPLUSB11 SFQOUTMINUSB11 WEIGHTLB11 WEIGHTRB11
XB11 SYNAPSEfastest SYNB11 0 DOUT13 WEIGHTLB11 WEIGHTRB11 INITIALB11
#lB111 SFQOUTPLUSB11 0 1p
#lB112 SFQOUTMINUSB11 0 1p

#ACTIVATION
XACT11 COMP5 XIN1 DOUT11 A4 DCIN DC4 DOUTL11 0  0 DOUTR12  0 DOUTL13 OUTPUT1GND OUTPUT1 OUTPUT2GND OUTPUT2   THRESH

#AXON FOR OUTPUT
XTRANSMIT1 TRANSMIT DOUTL11 XIN2 B4 A4 A6 DC4 DC6 DCCIN DCC4 OUTPUTAXON

#DELAYS
XDELAYACT1 DELAY10 DOUTR12 B4 B5 A6 A7 DC6 DC7  DELAYOUT1 0  DELAYOUT2 0
XDELAYTARGET DELAY14 ADJUSTTARGET1 B5 B6 A7 A8 DC7 DC8  DELAYOUTTARGET1  0 DELAYOUTTARGET2 0
#XDELAYTARGET2 DELAY103 ADJUSTTARGET2 B7 B8 A9 A10 DC9 DC10  DELAYOUTTARGET3 DELAYOUTTARGET3GND   DELAYOUTTARGET4 DELAYOUTTARGET4GND DELAYOUTTARGET5  DELAYOUTTARGET5GND 
XDELAYTARGET2 DELAY163 ADJUSTTARGET2 B7 B8 A9 A10 DC9 DC10  DELAYOUTTARGET3 DELAYOUTTARGET3GND   DELAYOUTTARGET4 DELAYOUTTARGET4GND DELAYOUTTARGET5  DELAYOUTTARGET5GND 


#LEARNING ALGORITHMS
#ASSUME DOUTFINAL1 0 DOUTFINAL2 0  DOUTFINAL3 0  0 DOUTFINAL4
#XMLP MLPNEW B6 B7 A8 A9 DELAYOUT1 DELAYOUT2 DELAYOUTTARGET1 DELAYOUTTARGET2 ACTNEXT1 ACTNEXT2 DC8 DC9 OUTPUTTARGET1L 0 OUTPUTTARGET2L 0 OUTPUTTARGET3L 0
#XDELAYTARGET2 DELAY18 ADJUSTTARGET2 B7 B8 A9 A10 DC9 dc10  DELAYOUTTARGET3GND DELAYOUTTARGET3  DELAYOUTTARGET4 DELAYOUTTARGET4GND  DELAYOUTTARGET5GND DELAYOUTTARGET5 
XMLP MLPNEW B6 B7 A8 A9 DELAYOUT1 DELAYOUT2 DELAYOUTTARGET1 DELAYOUTTARGET2 ACTNEXT1 ACTNEXT2 DC8 DC9  OUTPUTTARGET1L 0 OUTPUTTARGET2L 0 OUTPUTTARGET3L 0

XDELAYINPUT1 DELAY18 ADJUST11  B8  B9  A10 A11 DC10 DC11 DELAYOUTINPUT111 0 DELAYOUTINPUT112 0 DELAYOUTINPUT113 0 DELAYOUTINPUT114 0 DELAYOUTINPUT115 0 DELAYOUTINPUT116 0
XDELAYINPUT2 DELAY18 ADJUST12  B9  B10  A11 A12 DC11 DC12 DELAYOUTINPUT121 0 DELAYOUTINPUT122 0 DELAYOUTINPUT123 0 DELAYOUTINPUT124 0 DELAYOUTINPUT125 0 DELAYOUTINPUT126 0
XDELAYINPUTB1 DELAY18 ADJUSTB11  B10  B11  A12 A13 DC12 DC13 DELAYOUTINPUT1B1 0 DELAYOUTINPUT1B2 0 DELAYOUTINPUT1B3 0 DELAYOUTINPUT1B4 0 DELAYOUTINPUT1B5 0 DELAYOUTINPUT1B6 0

XDELAYact2 DELAY15 DOUTL13  B11 B12  A13 A14 DC13 DC14  DELAYOUTact111 0 0  DELAYOUTact112 DELAYOUTact113 0 0  DELAYOUTact114   DELAYOUTact115  0 0  DELAYOUTact116 


XPERCEPTRON11 PERCEPTRON  B13 B12  A14 A15  DELAYOUTINPUT111 DELAYOUTact111 DELAYOUTact112 OUTPUTTARGET1L DC15 DC14 INCR11 DECR11
XPERCEPTRON12 PERCEPTRON  B14 B13  A15 A16  DELAYOUTINPUT121 DELAYOUTact113 DELAYOUTact114 OUTPUTTARGET2L DC16 DC15 INCR12 DECR12
XPERCEPTRONB11 PERCEPTRON  XOUT2 B14  A16 A17  DELAYOUTINPUT1B1 DELAYOUTact115 DELAYOUTact116 OUTPUTTARGET3L DCOUT DC16 INCRB11 DECRB11

XCONV11 CONV A17 A18 DCC5 DCC4 INCR11 DECR11 SFQOUTPLUS11 SFQOUTMINUS11
XCONV12 CONV A18 A19 DCC6 DCC5 INCR12 DECR12 SFQOUTPLUS12 SFQOUTMINUS12
XCONVB11 CONV A19 XOUT1 DCCOUT DCC6 INCRB11 DECRB11 SFQOUTPLUSB11 SFQOUTMINUSB11

.ENDS 3NEURON2


.SUBCKT MLPNEW XIN1 XOUT1 XIN2 XOUT2 OI1 OI2 T1 T2 OJ1 OJ2 DCIN DCOUT OUTPUTTARGET1L OUTPUTTARGET1R OUTPUTTARGET2L OUTPUTTARGET2R OUTPUTTARGET3L OUTPUTTARGET3R
#Oi.T
Xand1  AND  B7 XIN1  XIN2 A9  OI1 T1 DC9 DCIN  andout1
#Oi.!Oj
Xand2  AND B8 B7 A9 A10 OI2 OJ1 DC10 DC9 andout2
#T.!Oj
Xand3  AND B9 B8 A10 A11 T2 OJ2 DC11 DC10 andout3
#D=Oi.T + Oi.!Oj + T.!Oj 
X3OR OR3 B9 XOUT1 XOUT2 A11   ANDOUT1 ANDOUT2 ANDOUT3 DCOUT DC11  OUTPUTTARGET1L OUTPUTTARGET1R OUTPUTTARGET2L OUTPUTTARGET2R OUTPUTTARGET3L OUTPUTTARGET3R 
.ENDS MLPNEW













.SUBCKT DELAY10 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 XOUT1  DC15 DC14      DELAYOUT9 0
XDELAY10 bfrsplit2 XOUT2 DELAYOUT9 A10   DC15 DCOUT      OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R
.ends DELAY10


.SUBCKT DELAY103 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R  OUTPUT3L OUTPUT3R

XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR XOUT2 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 bfrsplit3 XOUT1 DELAYOUT6 B7  DCOUT DC12 OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R

.ends DELAY103


.SUBCKT DELAY11 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR XOUT2 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 bfrsplit2 XOUT1 DELAYOUT10 B9   DCOUT DC16   OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R

.ends DELAY11




.SUBCKT DELAY14 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R

XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR A11 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 BFR B10 DELAYOUT10 B9   DC17 DC16   DELAYOUT11 0
XDELAY12 BFR A11 DELAYOUT11 A12   DC17 DC18  DELAYOUT12 0
XDELAY13 BFR B10 DELAYOUT12 XOUT1  DC19 DC18  DELAYOUT13 0
XDELAY14 bfrsplit2 XOUT2 DELAYOUT13 A12  DC19 DCOUT  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R
#XDELAY14 bfrsplit5 XOUT2 DELAYOUT13 A12  DC19 DCOUT  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R OUTPUT4L OUTPUT4R OUTPUT5L OUTPUT5R

.ends DELAY14


.SUBCKT DELAY143 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R

XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR A11 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 BFR B10 DELAYOUT10 B9   DC17 DC16   DELAYOUT11 0
XDELAY12 BFR A11 DELAYOUT11 A12   DC17 DC18  DELAYOUT12 0
XDELAY13 BFR B10 DELAYOUT12 XOUT1  DC19 DC18  DELAYOUT13 0
XDELAY14 bfrsplit3 XOUT2 DELAYOUT13 A12  DC19 DCOUT  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R
#XDELAY14 bfrsplit5 XOUT2 DELAYOUT13 A12  DC19 DCOUT  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R OUTPUT4L OUTPUT4R OUTPUT5L OUTPUT5R

.ends DELAY143

.SUBCKT DELAY15 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R OUTPUT4L OUTPUT4R OUTPUT5L OUTPUT5R OUTPUT6L OUTPUT6R
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR A11 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 BFR B10 DELAYOUT10 B9   DC17 DC16   DELAYOUT11 0
XDELAY12 BFR A11 DELAYOUT11 A12   DC17 DC18  DELAYOUT12 0
XDELAY13 BFR B10 DELAYOUT12 B11  DC19 DC18  DELAYOUT13 0
XDELAY14 BFR XOUT2 DELAYOUT13 A12  DC19 DC20  DELAYOUT14 0

XDELAY15 bfrsplit6 XOUT1 DELAYOUT14 B11 DCOUT DC20  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R OUTPUT4L OUTPUT4R OUTPUT5L OUTPUT5R OUTPUT6L OUTPUT6R

.ends DELAY15

.SUBCKT DELAY153 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R 
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR A11 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 BFR B10 DELAYOUT10 B9   DC17 DC16   DELAYOUT11 0
XDELAY12 BFR A11 DELAYOUT11 A12   DC17 DC18  DELAYOUT12 0
XDELAY13 BFR B10 DELAYOUT12 B11  DC19 DC18  DELAYOUT13 0
XDELAY14 BFR XOUT2 DELAYOUT13 A12  DC19 DC20  DELAYOUT14 0

XDELAY15 bfrsplit3 XOUT1 DELAYOUT14 B11 DCOUT DC20  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R 

.ends DELAY153



.SUBCKT DELAY16 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR A11 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 BFR B10 DELAYOUT10 B9   DC17 DC16   DELAYOUT11 0
XDELAY12 BFR A11 DELAYOUT11 A12   DC17 DC18  DELAYOUT12 0
XDELAY13 BFR B10 DELAYOUT12 B11  DC19 DC18  DELAYOUT13 0
XDELAY14 BFR A13 DELAYOUT13 A12  DC19 DC20  DELAYOUT14 0
XDELAY15 BFR XOUT1 DELAYOUT14 B11  DC21 DC20  DELAYOUT15 0
XDELAY16 bfrsplit2 A13 DELAYOUT15 XOUT2  DC21 DCOUT  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R
.ends DELAY16

.SUBCKT DELAY163 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR A11 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 BFR B10 DELAYOUT10 B9   DC17 DC16   DELAYOUT11 0
XDELAY12 BFR A11 DELAYOUT11 A12   DC17 DC18  DELAYOUT12 0
XDELAY13 BFR B10 DELAYOUT12 B11  DC19 DC18  DELAYOUT13 0
XDELAY14 BFR A13 DELAYOUT13 A12  DC19 DC20  DELAYOUT14 0
XDELAY15 BFR XOUT1 DELAYOUT14 B11  DC21 DC20  DELAYOUT15 0
XDELAY16 bfrsplit3 A13 DELAYOUT15 XOUT2  DC21 DCOUT  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R
.ends DELAY163


.SUBCKT DELAY18 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR A11 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 BFR B10 DELAYOUT10 B9   DC17 DC16   DELAYOUT11 0
XDELAY12 BFR A11 DELAYOUT11 A12   DC17 DC18  DELAYOUT12 0
XDELAY13 BFR B10 DELAYOUT12 B11  DC19 DC18  DELAYOUT13 0
XDELAY14 BFR A13 DELAYOUT13 A12  DC19 DC20  DELAYOUT14 0
XDELAY15 BFR B12 DELAYOUT14 B11  DC21 DC20  DELAYOUT15 0
XDELAY16 BFR A13 DELAYOUT15 A14  DC21 DC22  DELAYOUT16 0
XDELAY17 BFR B12 DELAYOUT16 XOUT1  DC23 DC22  DELAYOUT17 0
XDELAY18 bfrsplit3 XOUT2 DELAYOUT17 A14 DC23 DCOUT  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R  OUTPUT3L OUTPUT3R


.ends DELAY18

***    INPUTS  ***
IIN1 0 IN1 PWL(0 0 20P 0 1.55000e-09 0.00000e+00 1.55500e-09 2.00000e-03 1.60500e-09 2.00000e-03
+ 1.61000e-09 0.00000e+00 3.55000e-09 0.00000e+00 3.55500e-09 2.00000e-03
+ 3.60500e-09 2.00000e-03 3.61000e-09 0.00000e+00 5.55000e-09 0.00000e+00
+ 5.55500e-09 2.00000e-03 5.60500e-09 2.00000e-03 5.61000e-09 0.00000e+00
+ 7.55000e-09 0.00000e+00 7.55500e-09 2.00000e-03 7.60500e-09 2.00000e-03
+ 7.61000e-09 0.00000e+00 9.55000e-09 0.00000e+00 9.55500e-09 2.00000e-03
+ 9.60500e-09 2.00000e-03 9.61000e-09 0.00000e+00 1.15500e-08 0.00000e+00
+ 1.15550e-08 2.00000e-03 1.16050e-08 2.00000e-03 1.16100e-08 0.00000e+00
+ 1.35500e-08 0.00000e+00 1.35550e-08 2.00000e-03 1.36050e-08 2.00000e-03
+ 1.36100e-08 0.00000e+00 1.55500e-08 0.00000e+00 1.55550e-08 2.00000e-03
+ 1.56050e-08 2.00000e-03 1.56100e-08 0.00000e+00 1.75500e-08 0.00000e+00
+ 1.75550e-08 2.00000e-03 1.76050e-08 2.00000e-03 1.76100e-08 0.00000e+00
+ 1.95500e-08 0.00000e+00 1.95550e-08 2.00000e-03 1.96050e-08 2.00000e-03
+ 1.96100e-08 0.00000e+00 2.15500e-08 0.00000e+00 2.15550e-08 2.00000e-03
+ 2.16050e-08 2.00000e-03 2.16100e-08 0.00000e+00 2.35500e-08 0.00000e+00
+ 2.35550e-08 2.00000e-03 2.36050e-08 2.00000e-03 2.36100e-08 0.00000e+00
+ 2.55500e-08 0.00000e+00 2.55550e-08 2.00000e-03 2.56050e-08 2.00000e-03
+ 2.56100e-08 0.00000e+00 2.75500e-08 0.00000e+00 2.75550e-08 2.00000e-03
+ 2.76050e-08 2.00000e-03 2.76100e-08 0.00000e+00 2.95500e-08 0.00000e+00
+ 2.95550e-08 2.00000e-03 2.96050e-08 2.00000e-03 2.96100e-08 0.00000e+00
+ 3.15500e-08 0.00000e+00 3.15550e-08 2.00000e-03 3.16050e-08 2.00000e-03
+ 3.16100e-08 0.00000e+00 3.35500e-08 0.00000e+00 3.35550e-08 2.00000e-03
+ 3.36050e-08 2.00000e-03 3.36100e-08 0.00000e+00 3.55500e-08 0.00000e+00
+ 3.55550e-08 2.00000e-03 3.56050e-08 2.00000e-03 3.56100e-08 0.00000e+00
+ 3.75500e-08 0.00000e+00 3.75550e-08 2.00000e-03 3.76050e-08 2.00000e-03
+ 3.76100e-08 0.00000e+00 3.95500e-08 0.00000e+00 3.95550e-08 2.00000e-03
+ 3.96050e-08 2.00000e-03 3.96100e-08 0.00000e+00 4.15500e-08 0.00000e+00
+ 4.15550e-08 2.00000e-03 4.16050e-08 2.00000e-03 4.16100e-08 0.00000e+00
+ 4.35500e-08 0.00000e+00 4.35550e-08 2.00000e-03 4.36050e-08 2.00000e-03
+ 4.36100e-08 0.00000e+00 4.55500e-08 0.00000e+00 4.55550e-08 2.00000e-03
+ 4.56050e-08 2.00000e-03 4.56100e-08 0.00000e+00 4.75500e-08 0.00000e+00
+ 4.75550e-08 2.00000e-03 4.76050e-08 2.00000e-03 4.76100e-08 0.00000e+00
+ 4.95500e-08 0.00000e+00 4.95550e-08 2.00000e-03 4.96050e-08 2.00000e-03
+ 4.96100e-08 0.00000e+00 5.15500e-08 0.00000e+00 5.15550e-08 2.00000e-03
+ 5.16050e-08 2.00000e-03 5.16100e-08 0.00000e+00 5.35500e-08 0.00000e+00
+ 5.35550e-08 2.00000e-03 5.36050e-08 2.00000e-03 5.36100e-08 0.00000e+00
+ 5.55500e-08 0.00000e+00 5.55550e-08 2.00000e-03 5.56050e-08 2.00000e-03
+ 5.56100e-08 0.00000e+00 5.75500e-08 0.00000e+00 5.75550e-08 2.00000e-03
+ 5.76050e-08 2.00000e-03 5.76100e-08 0.00000e+00 5.95500e-08 0.00000e+00
+ 5.95550e-08 2.00000e-03 5.96050e-08 2.00000e-03 5.96100e-08 0.00000e+00
+ 6.15500e-08 0.00000e+00 6.15550e-08 2.00000e-03 6.16050e-08 2.00000e-03
+ 6.16100e-08 0.00000e+00 6.35500e-08 0.00000e+00 6.35550e-08 2.00000e-03
+ 6.36050e-08 2.00000e-03 6.36100e-08 0.00000e+00 6.55500e-08 0.00000e+00
+ 6.55550e-08 2.00000e-03 6.56050e-08 2.00000e-03 6.56100e-08 0.00000e+00
+ 6.75500e-08 0.00000e+00 6.75550e-08 2.00000e-03 6.76050e-08 2.00000e-03
+ 6.76100e-08 0.00000e+00 6.95500e-08 0.00000e+00 6.95550e-08 2.00000e-03
+ 6.96050e-08 2.00000e-03 6.96100e-08 0.00000e+00 7.15500e-08 0.00000e+00
+ 7.15550e-08 2.00000e-03 7.16050e-08 2.00000e-03 7.16100e-08 0.00000e+00
+ 7.35500e-08 0.00000e+00 7.35550e-08 2.00000e-03 7.36050e-08 2.00000e-03
+ 7.36100e-08 0.00000e+00 7.55500e-08 0.00000e+00 7.55550e-08 2.00000e-03
+ 7.56050e-08 2.00000e-03 7.56100e-08 0.00000e+00 7.75500e-08 0.00000e+00
+ 7.75550e-08 2.00000e-03 7.76050e-08 2.00000e-03 7.76100e-08 0.00000e+00
+ 7.95500e-08 0.00000e+00 7.95550e-08 2.00000e-03 7.96050e-08 2.00000e-03
+ 7.96100e-08 0.00000e+00 8.15500e-08 0.00000e+00 8.15550e-08 2.00000e-03
+ 8.16050e-08 2.00000e-03 8.16100e-08 0.00000e+00 8.35500e-08 0.00000e+00
+ 8.35550e-08 2.00000e-03 8.36050e-08 2.00000e-03 8.36100e-08 0.00000e+00
+ 8.55500e-08 0.00000e+00 8.55550e-08 2.00000e-03 8.56050e-08 2.00000e-03
+ 8.56100e-08 0.00000e+00 8.75500e-08 0.00000e+00 8.75550e-08 2.00000e-03
+ 8.76050e-08 2.00000e-03 8.76100e-08 0.00000e+00 8.95500e-08 0.00000e+00
+ 8.95550e-08 2.00000e-03 8.96050e-08 2.00000e-03 8.96100e-08 0.00000e+00
+ 9.15500e-08 0.00000e+00 9.15550e-08 2.00000e-03 9.16050e-08 2.00000e-03
+ 9.16100e-08 0.00000e+00 9.35500e-08 0.00000e+00 9.35550e-08 2.00000e-03
+ 9.36050e-08 2.00000e-03 9.36100e-08 0.00000e+00 9.55500e-08 0.00000e+00
+ 9.55550e-08 2.00000e-03 9.56050e-08 2.00000e-03 9.56100e-08 0.00000e+00
+ 9.75500e-08 0.00000e+00 9.75550e-08 2.00000e-03 9.76050e-08 2.00000e-03
+ 9.76100e-08 0.00000e+00 9.95500e-08 0.00000e+00 9.95550e-08 2.00000e-03
+ 9.96050e-08 2.00000e-03 9.96100e-08 0.00000e+00 1.01550e-07 0.00000e+00
+ 1.01555e-07 2.00000e-03 1.01605e-07 2.00000e-03 1.01610e-07 0.00000e+00
+ 1.03550e-07 0.00000e+00 1.03555e-07 2.00000e-03 1.03605e-07 2.00000e-03
+ 1.03610e-07 0.00000e+00 1.05550e-07 0.00000e+00 1.05555e-07 2.00000e-03
+ 1.05605e-07 2.00000e-03 1.05610e-07 0.00000e+00 1.07550e-07 0.00000e+00
+ 1.07555e-07 2.00000e-03 1.07605e-07 2.00000e-03 1.07610e-07 0.00000e+00
+ 1.09550e-07 0.00000e+00 1.09555e-07 2.00000e-03 1.09605e-07 2.00000e-03
+ 1.09610e-07 0.00000e+00 1.11550e-07 0.00000e+00 1.11555e-07 2.00000e-03
+ 1.11605e-07 2.00000e-03 1.11610e-07 0.00000e+00 1.13550e-07 0.00000e+00
+ 1.13555e-07 2.00000e-03 1.13605e-07 2.00000e-03 1.13610e-07 0.00000e+00
+ 1.15550e-07 0.00000e+00 1.15555e-07 2.00000e-03 1.15605e-07 2.00000e-03
+ 1.15610e-07 0.00000e+00 1.17550e-07 0.00000e+00 1.17555e-07 2.00000e-03
+ 1.17605e-07 2.00000e-03 1.17610e-07 0.00000e+00 1.19550e-07 0.00000e+00
+ 1.19555e-07 2.00000e-03 1.19605e-07 2.00000e-03 1.19610e-07 0.00000e+00)
IIN2 0 IN2 PWL(0 0 20P 0 2.55000e-09 0.00000e+00 2.55500e-09 2.00000e-03 2.60500e-09 2.00000e-03
+ 2.61000e-09 0.00000e+00 3.55000e-09 0.00000e+00 3.55500e-09 2.00000e-03
+ 3.60500e-09 2.00000e-03 3.61000e-09 0.00000e+00 6.55000e-09 0.00000e+00
+ 6.55500e-09 2.00000e-03 6.60500e-09 2.00000e-03 6.61000e-09 0.00000e+00
+ 7.55000e-09 0.00000e+00 7.55500e-09 2.00000e-03 7.60500e-09 2.00000e-03
+ 7.61000e-09 0.00000e+00 1.05500e-08 0.00000e+00 1.05550e-08 2.00000e-03
+ 1.06050e-08 2.00000e-03 1.06100e-08 0.00000e+00 1.15500e-08 0.00000e+00
+ 1.15550e-08 2.00000e-03 1.16050e-08 2.00000e-03 1.16100e-08 0.00000e+00
+ 1.45500e-08 0.00000e+00 1.45550e-08 2.00000e-03 1.46050e-08 2.00000e-03
+ 1.46100e-08 0.00000e+00 1.55500e-08 0.00000e+00 1.55550e-08 2.00000e-03
+ 1.56050e-08 2.00000e-03 1.56100e-08 0.00000e+00 1.85500e-08 0.00000e+00
+ 1.85550e-08 2.00000e-03 1.86050e-08 2.00000e-03 1.86100e-08 0.00000e+00
+ 1.95500e-08 0.00000e+00 1.95550e-08 2.00000e-03 1.96050e-08 2.00000e-03
+ 1.96100e-08 0.00000e+00 2.25500e-08 0.00000e+00 2.25550e-08 2.00000e-03
+ 2.26050e-08 2.00000e-03 2.26100e-08 0.00000e+00 2.35500e-08 0.00000e+00
+ 2.35550e-08 2.00000e-03 2.36050e-08 2.00000e-03 2.36100e-08 0.00000e+00
+ 2.65500e-08 0.00000e+00 2.65550e-08 2.00000e-03 2.66050e-08 2.00000e-03
+ 2.66100e-08 0.00000e+00 2.75500e-08 0.00000e+00 2.75550e-08 2.00000e-03
+ 2.76050e-08 2.00000e-03 2.76100e-08 0.00000e+00 3.05500e-08 0.00000e+00
+ 3.05550e-08 2.00000e-03 3.06050e-08 2.00000e-03 3.06100e-08 0.00000e+00
+ 3.15500e-08 0.00000e+00 3.15550e-08 2.00000e-03 3.16050e-08 2.00000e-03
+ 3.16100e-08 0.00000e+00 3.45500e-08 0.00000e+00 3.45550e-08 2.00000e-03
+ 3.46050e-08 2.00000e-03 3.46100e-08 0.00000e+00 3.55500e-08 0.00000e+00
+ 3.55550e-08 2.00000e-03 3.56050e-08 2.00000e-03 3.56100e-08 0.00000e+00
+ 3.85500e-08 0.00000e+00 3.85550e-08 2.00000e-03 3.86050e-08 2.00000e-03
+ 3.86100e-08 0.00000e+00 3.95500e-08 0.00000e+00 3.95550e-08 2.00000e-03
+ 3.96050e-08 2.00000e-03 3.96100e-08 0.00000e+00 4.25500e-08 0.00000e+00
+ 4.25550e-08 2.00000e-03 4.26050e-08 2.00000e-03 4.26100e-08 0.00000e+00
+ 4.35500e-08 0.00000e+00 4.35550e-08 2.00000e-03 4.36050e-08 2.00000e-03
+ 4.36100e-08 0.00000e+00 4.65500e-08 0.00000e+00 4.65550e-08 2.00000e-03
+ 4.66050e-08 2.00000e-03 4.66100e-08 0.00000e+00 4.75500e-08 0.00000e+00
+ 4.75550e-08 2.00000e-03 4.76050e-08 2.00000e-03 4.76100e-08 0.00000e+00
+ 5.05500e-08 0.00000e+00 5.05550e-08 2.00000e-03 5.06050e-08 2.00000e-03
+ 5.06100e-08 0.00000e+00 5.15500e-08 0.00000e+00 5.15550e-08 2.00000e-03
+ 5.16050e-08 2.00000e-03 5.16100e-08 0.00000e+00 5.45500e-08 0.00000e+00
+ 5.45550e-08 2.00000e-03 5.46050e-08 2.00000e-03 5.46100e-08 0.00000e+00
+ 5.55500e-08 0.00000e+00 5.55550e-08 2.00000e-03 5.56050e-08 2.00000e-03
+ 5.56100e-08 0.00000e+00 5.85500e-08 0.00000e+00 5.85550e-08 2.00000e-03
+ 5.86050e-08 2.00000e-03 5.86100e-08 0.00000e+00 5.95500e-08 0.00000e+00
+ 5.95550e-08 2.00000e-03 5.96050e-08 2.00000e-03 5.96100e-08 0.00000e+00
+ 6.25500e-08 0.00000e+00 6.25550e-08 2.00000e-03 6.26050e-08 2.00000e-03
+ 6.26100e-08 0.00000e+00 6.35500e-08 0.00000e+00 6.35550e-08 2.00000e-03
+ 6.36050e-08 2.00000e-03 6.36100e-08 0.00000e+00 6.65500e-08 0.00000e+00
+ 6.65550e-08 2.00000e-03 6.66050e-08 2.00000e-03 6.66100e-08 0.00000e+00
+ 6.75500e-08 0.00000e+00 6.75550e-08 2.00000e-03 6.76050e-08 2.00000e-03
+ 6.76100e-08 0.00000e+00 7.05500e-08 0.00000e+00 7.05550e-08 2.00000e-03
+ 7.06050e-08 2.00000e-03 7.06100e-08 0.00000e+00 7.15500e-08 0.00000e+00
+ 7.15550e-08 2.00000e-03 7.16050e-08 2.00000e-03 7.16100e-08 0.00000e+00
+ 7.45500e-08 0.00000e+00 7.45550e-08 2.00000e-03 7.46050e-08 2.00000e-03
+ 7.46100e-08 0.00000e+00 7.55500e-08 0.00000e+00 7.55550e-08 2.00000e-03
+ 7.56050e-08 2.00000e-03 7.56100e-08 0.00000e+00 7.85500e-08 0.00000e+00
+ 7.85550e-08 2.00000e-03 7.86050e-08 2.00000e-03 7.86100e-08 0.00000e+00
+ 7.95500e-08 0.00000e+00 7.95550e-08 2.00000e-03 7.96050e-08 2.00000e-03
+ 7.96100e-08 0.00000e+00 8.25500e-08 0.00000e+00 8.25550e-08 2.00000e-03
+ 8.26050e-08 2.00000e-03 8.26100e-08 0.00000e+00 8.35500e-08 0.00000e+00
+ 8.35550e-08 2.00000e-03 8.36050e-08 2.00000e-03 8.36100e-08 0.00000e+00
+ 8.65500e-08 0.00000e+00 8.65550e-08 2.00000e-03 8.66050e-08 2.00000e-03
+ 8.66100e-08 0.00000e+00 8.75500e-08 0.00000e+00 8.75550e-08 2.00000e-03
+ 8.76050e-08 2.00000e-03 8.76100e-08 0.00000e+00 9.05500e-08 0.00000e+00
+ 9.05550e-08 2.00000e-03 9.06050e-08 2.00000e-03 9.06100e-08 0.00000e+00
+ 9.15500e-08 0.00000e+00 9.15550e-08 2.00000e-03 9.16050e-08 2.00000e-03
+ 9.16100e-08 0.00000e+00 9.45500e-08 0.00000e+00 9.45550e-08 2.00000e-03
+ 9.46050e-08 2.00000e-03 9.46100e-08 0.00000e+00 9.55500e-08 0.00000e+00
+ 9.55550e-08 2.00000e-03 9.56050e-08 2.00000e-03 9.56100e-08 0.00000e+00
+ 9.85500e-08 0.00000e+00 9.85550e-08 2.00000e-03 9.86050e-08 2.00000e-03
+ 9.86100e-08 0.00000e+00 9.95500e-08 0.00000e+00 9.95550e-08 2.00000e-03
+ 9.96050e-08 2.00000e-03 9.96100e-08 0.00000e+00 1.02550e-07 0.00000e+00
+ 1.02555e-07 2.00000e-03 1.02605e-07 2.00000e-03 1.02610e-07 0.00000e+00
+ 1.03550e-07 0.00000e+00 1.03555e-07 2.00000e-03 1.03605e-07 2.00000e-03
+ 1.03610e-07 0.00000e+00 1.06550e-07 0.00000e+00 1.06555e-07 2.00000e-03
+ 1.06605e-07 2.00000e-03 1.06610e-07 0.00000e+00 1.07550e-07 0.00000e+00
+ 1.07555e-07 2.00000e-03 1.07605e-07 2.00000e-03 1.07610e-07 0.00000e+00
+ 1.10550e-07 0.00000e+00 1.10555e-07 2.00000e-03 1.10605e-07 2.00000e-03
+ 1.10610e-07 0.00000e+00 1.11550e-07 0.00000e+00 1.11555e-07 2.00000e-03
+ 1.11605e-07 2.00000e-03 1.11610e-07 0.00000e+00 1.14550e-07 0.00000e+00
+ 1.14555e-07 2.00000e-03 1.14605e-07 2.00000e-03 1.14610e-07 0.00000e+00
+ 1.15550e-07 0.00000e+00 1.15555e-07 2.00000e-03 1.15605e-07 2.00000e-03
+ 1.15610e-07 0.00000e+00 1.18550e-07 0.00000e+00 1.18555e-07 2.00000e-03
+ 1.18605e-07 2.00000e-03 1.18610e-07 0.00000e+00 1.19550e-07 0.00000e+00
+ 1.19555e-07 2.00000e-03 1.19605e-07 2.00000e-03 1.19610e-07 0.00000e+00)
IINBIAS1 0 INB11 pulse(0 0.002 550p 5p 5p 50p 1000p)
ITARGET 0 TARGET0  PWL(0 0 20P 0 3.55000e-09 0.00000e+00 3.55500e-09 2.00000e-03 3.60500e-09 2.00000e-03
+ 3.61000e-09 0.00000e+00 7.55000e-09 0.00000e+00 7.55500e-09 2.00000e-03
+ 7.60500e-09 2.00000e-03 7.61000e-09 0.00000e+00 1.15500e-08 0.00000e+00
+ 1.15550e-08 2.00000e-03 1.16050e-08 2.00000e-03 1.16100e-08 0.00000e+00
+ 1.55500e-08 0.00000e+00 1.55550e-08 2.00000e-03 1.56050e-08 2.00000e-03
+ 1.56100e-08 0.00000e+00 1.95500e-08 0.00000e+00 1.95550e-08 2.00000e-03
+ 1.96050e-08 2.00000e-03 1.96100e-08 0.00000e+00 2.35500e-08 0.00000e+00
+ 2.35550e-08 2.00000e-03 2.36050e-08 2.00000e-03 2.36100e-08 0.00000e+00
+ 2.75500e-08 0.00000e+00 2.75550e-08 2.00000e-03 2.76050e-08 2.00000e-03
+ 2.76100e-08 0.00000e+00 3.15500e-08 0.00000e+00 3.15550e-08 2.00000e-03
+ 3.16050e-08 2.00000e-03 3.16100e-08 0.00000e+00 3.55500e-08 0.00000e+00
+ 3.55550e-08 2.00000e-03 3.56050e-08 2.00000e-03 3.56100e-08 0.00000e+00
+ 3.95500e-08 0.00000e+00 3.95550e-08 2.00000e-03 3.96050e-08 2.00000e-03
+ 3.96100e-08 0.00000e+00 4.35500e-08 0.00000e+00 4.35550e-08 2.00000e-03
+ 4.36050e-08 2.00000e-03 4.36100e-08 0.00000e+00 4.75500e-08 0.00000e+00
+ 4.75550e-08 2.00000e-03 4.76050e-08 2.00000e-03 4.76100e-08 0.00000e+00
+ 5.15500e-08 0.00000e+00 5.15550e-08 2.00000e-03 5.16050e-08 2.00000e-03
+ 5.16100e-08 0.00000e+00 5.55500e-08 0.00000e+00 5.55550e-08 2.00000e-03
+ 5.56050e-08 2.00000e-03 5.56100e-08 0.00000e+00 5.95500e-08 0.00000e+00
+ 5.95550e-08 2.00000e-03 5.96050e-08 2.00000e-03 5.96100e-08 0.00000e+00
+ 6.35500e-08 0.00000e+00 6.35550e-08 2.00000e-03 6.36050e-08 2.00000e-03
+ 6.36100e-08 0.00000e+00 6.75500e-08 0.00000e+00 6.75550e-08 2.00000e-03
+ 6.76050e-08 2.00000e-03 6.76100e-08 0.00000e+00 7.15500e-08 0.00000e+00
+ 7.15550e-08 2.00000e-03 7.16050e-08 2.00000e-03 7.16100e-08 0.00000e+00
+ 7.55500e-08 0.00000e+00 7.55550e-08 2.00000e-03 7.56050e-08 2.00000e-03
+ 7.56100e-08 0.00000e+00 7.95500e-08 0.00000e+00 7.95550e-08 2.00000e-03
+ 7.96050e-08 2.00000e-03 7.96100e-08 0.00000e+00 8.35500e-08 0.00000e+00
+ 8.35550e-08 2.00000e-03 8.36050e-08 2.00000e-03 8.36100e-08 0.00000e+00
+ 8.75500e-08 0.00000e+00 8.75550e-08 2.00000e-03 8.76050e-08 2.00000e-03
+ 8.76100e-08 0.00000e+00 9.15500e-08 0.00000e+00 9.15550e-08 2.00000e-03
+ 9.16050e-08 2.00000e-03 9.16100e-08 0.00000e+00 9.55500e-08 0.00000e+00
+ 9.55550e-08 2.00000e-03 9.56050e-08 2.00000e-03 9.56100e-08 0.00000e+00
+ 9.95500e-08 0.00000e+00 9.95550e-08 2.00000e-03 9.96050e-08 2.00000e-03
+ 9.96100e-08 0.00000e+00 1.03550e-07 0.00000e+00 1.03555e-07 2.00000e-03
+ 1.03605e-07 2.00000e-03 1.03610e-07 0.00000e+00 1.07550e-07 0.00000e+00
+ 1.07555e-07 2.00000e-03 1.07605e-07 2.00000e-03 1.07610e-07 0.00000e+00
+ 1.11550e-07 0.00000e+00 1.11555e-07 2.00000e-03 1.11605e-07 2.00000e-03
+ 1.11610e-07 0.00000e+00 1.15550e-07 0.00000e+00 1.15555e-07 2.00000e-03
+ 1.15605e-07 2.00000e-03 1.15610e-07 0.00000e+00 1.19550e-07 0.00000e+00
+ 1.19555e-07 2.00000e-03 1.19605e-07 2.00000e-03 1.19610e-07 0.00000e+00)
Iactualsynbias21 0 ACTUALSYNB21x PWL(0 0 6.4000e-10 0.0000e+00 6.6500e-10 6.7000e-04 7.0000e-10 0.0000e+00
+ 8.4000e-10 0.0000e+00 8.6500e-10 6.7000e-04 9.0000e-10 0.0000e+00
+ 1.0400e-09 0.0000e+00 1.0650e-09 6.7000e-04 1.1000e-09 0.0000e+00
+ 1.2400e-09 0.0000e+00 1.2650e-09 6.7000e-04 1.3000e-09 0.0000e+00
+ 1.4400e-09 0.0000e+00 1.4650e-09 6.7000e-04 1.5000e-09 0.0000e+00
+ 1.6400e-09 0.0000e+00 1.6650e-09 6.7000e-04 1.7000e-09 0.0000e+00
+ 1.8400e-09 0.0000e+00 1.8650e-09 6.7000e-04 1.9000e-09 0.0000e+00
+ 2.0400e-09 0.0000e+00 2.0650e-09 6.7000e-04 2.1000e-09 0.0000e+00
+ 2.2400e-09 0.0000e+00 2.2650e-09 6.7000e-04 2.3000e-09 0.0000e+00
+ 2.4400e-09 0.0000e+00 2.4650e-09 6.7000e-04 2.5000e-09 0.0000e+00
+ 2.6400e-09 0.0000e+00 2.6650e-09 6.7000e-04 2.7000e-09 0.0000e+00
+ 2.8400e-09 0.0000e+00 2.8650e-09 6.7000e-04 2.9000e-09 0.0000e+00
+ 3.0400e-09 0.0000e+00 3.0650e-09 6.7000e-04 3.1000e-09 0.0000e+00
+ 3.2400e-09 0.0000e+00 3.2650e-09 6.7000e-04 3.3000e-09 0.0000e+00
+ 3.4400e-09 0.0000e+00 3.4650e-09 6.7000e-04 3.5000e-09 0.0000e+00
+ 3.6400e-09 0.0000e+00 3.6650e-09 6.7000e-04 3.7000e-09 0.0000e+00
+ 3.8400e-09 0.0000e+00 3.8650e-09 6.7000e-04 3.9000e-09 0.0000e+00
+ 4.0400e-09 0.0000e+00 4.0650e-09 6.7000e-04 4.1000e-09 0.0000e+00
+ 4.2400e-09 0.0000e+00 4.2650e-09 6.7000e-04 4.3000e-09 0.0000e+00
+ 4.4400e-09 0.0000e+00 4.4650e-09 6.7000e-04 4.5000e-09 0.0000e+00
+ 4.6400e-09 0.0000e+00 4.6650e-09 6.7000e-04 4.7000e-09 0.0000e+00
+ 4.8400e-09 0.0000e+00 4.8650e-09 6.7000e-04 4.9000e-09 0.0000e+00
+ 5.0400e-09 0.0000e+00 5.0650e-09 6.7000e-04 5.1000e-09 0.0000e+00
+ 5.2400e-09 0.0000e+00 5.2650e-09 6.7000e-04 5.3000e-09 0.0000e+00
+ 5.4400e-09 0.0000e+00 5.4650e-09 6.7000e-04 5.5000e-09 0.0000e+00
+ 5.6400e-09 0.0000e+00 5.6650e-09 6.7000e-04 5.7000e-09 0.0000e+00
+ 5.8400e-09 0.0000e+00 5.8650e-09 6.7000e-04 5.9000e-09 0.0000e+00
+ 6.0400e-09 0.0000e+00 6.0650e-09 6.7000e-04 6.1000e-09 0.0000e+00
+ 6.2400e-09 0.0000e+00 6.2650e-09 6.7000e-04 6.3000e-09 0.0000e+00
+ 6.4400e-09 0.0000e+00 6.4650e-09 6.7000e-04 6.5000e-09 0.0000e+00
+ 6.6400e-09 0.0000e+00 6.6650e-09 6.7000e-04 6.7000e-09 0.0000e+00
+ 6.8400e-09 0.0000e+00 6.8650e-09 6.7000e-04 6.9000e-09 0.0000e+00
+ 7.0400e-09 0.0000e+00 7.0650e-09 6.7000e-04 7.1000e-09 0.0000e+00
+ 7.2400e-09 0.0000e+00 7.2650e-09 6.7000e-04 7.3000e-09 0.0000e+00
+ 7.4400e-09 0.0000e+00 7.4650e-09 6.7000e-04 7.5000e-09 0.0000e+00
+ 7.6400e-09 0.0000e+00 7.6650e-09 6.7000e-04 7.7000e-09 0.0000e+00
+ 7.8400e-09 0.0000e+00 7.8650e-09 6.7000e-04 7.9000e-09 0.0000e+00
+ 8.0400e-09 0.0000e+00 8.0650e-09 6.7000e-04 8.1000e-09 0.0000e+00
+ 8.2400e-09 0.0000e+00 8.2650e-09 6.7000e-04 8.3000e-09 0.0000e+00
+ 8.4400e-09 0.0000e+00 8.4650e-09 6.7000e-04 8.5000e-09 0.0000e+00
+ 8.6400e-09 0.0000e+00 8.6650e-09 6.7000e-04 8.7000e-09 0.0000e+00
+ 8.8400e-09 0.0000e+00 8.8650e-09 6.7000e-04 8.9000e-09 0.0000e+00
+ 9.0400e-09 0.0000e+00 9.0650e-09 6.7000e-04 9.1000e-09 0.0000e+00
+ 9.2400e-09 0.0000e+00 9.2650e-09 6.7000e-04 9.3000e-09 0.0000e+00
+ 9.4400e-09 0.0000e+00 9.4650e-09 6.7000e-04 9.5000e-09 0.0000e+00
+ 9.6400e-09 0.0000e+00 9.6650e-09 6.7000e-04 9.7000e-09 0.0000e+00
+ 9.8400e-09 0.0000e+00 9.8650e-09 6.7000e-04 9.9000e-09 0.0000e+00
+ 1.0040e-08 0.0000e+00 1.0065e-08 6.7000e-04 1.0100e-08 0.0000e+00
+ 1.0240e-08 0.0000e+00 1.0265e-08 6.7000e-04 1.0300e-08 0.0000e+00
+ 1.0440e-08 0.0000e+00 1.0465e-08 6.7000e-04 1.0500e-08 0.0000e+00
+ 1.0640e-08 0.0000e+00 1.0665e-08 6.7000e-04 1.0700e-08 0.0000e+00
+ 1.0840e-08 0.0000e+00 1.0865e-08 6.7000e-04 1.0900e-08 0.0000e+00
+ 1.1040e-08 0.0000e+00 1.1065e-08 6.7000e-04 1.1100e-08 0.0000e+00
+ 1.1240e-08 0.0000e+00 1.1265e-08 6.7000e-04 1.1300e-08 0.0000e+00
+ 1.1440e-08 0.0000e+00 1.1465e-08 6.7000e-04 1.1500e-08 0.0000e+00
+ 1.1640e-08 0.0000e+00 1.1665e-08 6.7000e-04 1.1700e-08 0.0000e+00
+ 1.1840e-08 0.0000e+00 1.1865e-08 6.7000e-04 1.1900e-08 0.0000e+00
+ 1.2040e-08 0.0000e+00 1.2065e-08 6.7000e-04 1.2100e-08 0.0000e+00
+ 1.2240e-08 0.0000e+00 1.2265e-08 6.7000e-04 1.2300e-08 0.0000e+00
+ 1.2440e-08 0.0000e+00 1.2465e-08 6.7000e-04 1.2500e-08 0.0000e+00
+ 1.2640e-08 0.0000e+00 1.2665e-08 6.7000e-04 1.2700e-08 0.0000e+00
+ 1.2840e-08 0.0000e+00 1.2865e-08 6.7000e-04 1.2900e-08 0.0000e+00
+ 1.3040e-08 0.0000e+00 1.3065e-08 6.7000e-04 1.3100e-08 0.0000e+00
+ 1.3240e-08 0.0000e+00 1.3265e-08 6.7000e-04 1.3300e-08 0.0000e+00
+ 1.3440e-08 0.0000e+00 1.3465e-08 6.7000e-04 1.3500e-08 0.0000e+00
+ 1.3640e-08 0.0000e+00 1.3665e-08 6.7000e-04 1.3700e-08 0.0000e+00
+ 1.3840e-08 0.0000e+00 1.3865e-08 6.7000e-04 1.3900e-08 0.0000e+00
+ 1.4040e-08 0.0000e+00 1.4065e-08 6.7000e-04 1.4100e-08 0.0000e+00
+ 1.4240e-08 0.0000e+00 1.4265e-08 6.7000e-04 1.4300e-08 0.0000e+00
+ 1.4440e-08 0.0000e+00 1.4465e-08 6.7000e-04 1.4500e-08 0.0000e+00
+ 1.4640e-08 0.0000e+00 1.4665e-08 6.7000e-04 1.4700e-08 0.0000e+00
+ 1.4840e-08 0.0000e+00 1.4865e-08 6.7000e-04 1.4900e-08 0.0000e+00
+ 1.5040e-08 0.0000e+00 1.5065e-08 6.7000e-04 1.5100e-08 0.0000e+00
+ 1.5240e-08 0.0000e+00 1.5265e-08 6.7000e-04 1.5300e-08 0.0000e+00
+ 1.5440e-08 0.0000e+00 1.5465e-08 6.7000e-04 1.5500e-08 0.0000e+00
+ 1.5640e-08 0.0000e+00 1.5665e-08 6.7000e-04 1.5700e-08 0.0000e+00
+ 1.5840e-08 0.0000e+00 1.5865e-08 6.7000e-04 1.5900e-08 0.0000e+00
+ 1.6040e-08 0.0000e+00 1.6065e-08 6.7000e-04 1.6100e-08 0.0000e+00
+ 1.6240e-08 0.0000e+00 1.6265e-08 6.7000e-04 1.6300e-08 0.0000e+00
+ 1.6440e-08 0.0000e+00 1.6465e-08 6.7000e-04 1.6500e-08 0.0000e+00
+ 1.6640e-08 0.0000e+00 1.6665e-08 6.7000e-04 1.6700e-08 0.0000e+00
+ 1.6840e-08 0.0000e+00 1.6865e-08 6.7000e-04 1.6900e-08 0.0000e+00
+ 1.7040e-08 0.0000e+00 1.7065e-08 6.7000e-04 1.7100e-08 0.0000e+00
+ 1.7240e-08 0.0000e+00 1.7265e-08 6.7000e-04 1.7300e-08 0.0000e+00
+ 1.7440e-08 0.0000e+00 1.7465e-08 6.7000e-04 1.7500e-08 0.0000e+00
+ 1.7640e-08 0.0000e+00 1.7665e-08 6.7000e-04 1.7700e-08 0.0000e+00
+ 1.7840e-08 0.0000e+00 1.7865e-08 6.7000e-04 1.7900e-08 0.0000e+00
+ 1.8040e-08 0.0000e+00 1.8065e-08 6.7000e-04 1.8100e-08 0.0000e+00
+ 1.8240e-08 0.0000e+00 1.8265e-08 6.7000e-04 1.8300e-08 0.0000e+00
+ 1.8440e-08 0.0000e+00 1.8465e-08 6.7000e-04 1.8500e-08 0.0000e+00
+ 1.8640e-08 0.0000e+00 1.8665e-08 6.7000e-04 1.8700e-08 0.0000e+00
+ 1.8840e-08 0.0000e+00 1.8865e-08 6.7000e-04 1.8900e-08 0.0000e+00
+ 1.9040e-08 0.0000e+00 1.9065e-08 6.7000e-04 1.9100e-08 0.0000e+00
+ 1.9240e-08 0.0000e+00 1.9265e-08 6.7000e-04 1.9300e-08 0.0000e+00
+ 1.9440e-08 0.0000e+00 1.9465e-08 6.7000e-04 1.9500e-08 0.0000e+00
+ 1.9640e-08 0.0000e+00 1.9665e-08 6.7000e-04 1.9700e-08 0.0000e+00
+ 1.9840e-08 0.0000e+00 1.9865e-08 6.7000e-04 1.9900e-08 0.0000e+00
+ 2.0040e-08 0.0000e+00 2.0065e-08 6.7000e-04 2.0100e-08 0.0000e+00
+ 2.0240e-08 0.0000e+00 2.0265e-08 6.7000e-04 2.0300e-08 0.0000e+00
+ 2.0440e-08 0.0000e+00 2.0465e-08 6.7000e-04 2.0500e-08 0.0000e+00
+ 2.0640e-08 0.0000e+00 2.0665e-08 6.7000e-04 2.0700e-08 0.0000e+00
+ 2.0840e-08 0.0000e+00 2.0865e-08 6.7000e-04 2.0900e-08 0.0000e+00
+ 2.1040e-08 0.0000e+00 2.1065e-08 6.7000e-04 2.1100e-08 0.0000e+00
+ 2.1240e-08 0.0000e+00 2.1265e-08 6.7000e-04 2.1300e-08 0.0000e+00
+ 2.1440e-08 0.0000e+00 2.1465e-08 6.7000e-04 2.1500e-08 0.0000e+00
+ 2.1640e-08 0.0000e+00 2.1665e-08 6.7000e-04 2.1700e-08 0.0000e+00
+ 2.1840e-08 0.0000e+00 2.1865e-08 6.7000e-04 2.1900e-08 0.0000e+00
+ 2.2040e-08 0.0000e+00 2.2065e-08 6.7000e-04 2.2100e-08 0.0000e+00
+ 2.2240e-08 0.0000e+00 2.2265e-08 6.7000e-04 2.2300e-08 0.0000e+00
+ 2.2440e-08 0.0000e+00 2.2465e-08 6.7000e-04 2.2500e-08 0.0000e+00
+ 2.2640e-08 0.0000e+00 2.2665e-08 6.7000e-04 2.2700e-08 0.0000e+00
+ 2.2840e-08 0.0000e+00 2.2865e-08 6.7000e-04 2.2900e-08 0.0000e+00
+ 2.3040e-08 0.0000e+00 2.3065e-08 6.7000e-04 2.3100e-08 0.0000e+00
+ 2.3240e-08 0.0000e+00 2.3265e-08 6.7000e-04 2.3300e-08 0.0000e+00
+ 2.3440e-08 0.0000e+00 2.3465e-08 6.7000e-04 2.3500e-08 0.0000e+00
+ 2.3640e-08 0.0000e+00 2.3665e-08 6.7000e-04 2.3700e-08 0.0000e+00
+ 2.3840e-08 0.0000e+00 2.3865e-08 6.7000e-04 2.3900e-08 0.0000e+00
+ 2.4040e-08 0.0000e+00 2.4065e-08 6.7000e-04 2.4100e-08 0.0000e+00
+ 2.4240e-08 0.0000e+00 2.4265e-08 6.7000e-04 2.4300e-08 0.0000e+00
+ 2.4440e-08 0.0000e+00 2.4465e-08 6.7000e-04 2.4500e-08 0.0000e+00
+ 2.4640e-08 0.0000e+00 2.4665e-08 6.7000e-04 2.4700e-08 0.0000e+00
+ 2.4840e-08 0.0000e+00 2.4865e-08 6.7000e-04 2.4900e-08 0.0000e+00
+ 2.5040e-08 0.0000e+00 2.5065e-08 6.7000e-04 2.5100e-08 0.0000e+00
+ 2.5240e-08 0.0000e+00 2.5265e-08 6.7000e-04 2.5300e-08 0.0000e+00
+ 2.5440e-08 0.0000e+00 2.5465e-08 6.7000e-04 2.5500e-08 0.0000e+00
+ 2.5640e-08 0.0000e+00 2.5665e-08 6.7000e-04 2.5700e-08 0.0000e+00
+ 2.5840e-08 0.0000e+00 2.5865e-08 6.7000e-04 2.5900e-08 0.0000e+00
+ 2.6040e-08 0.0000e+00 2.6065e-08 6.7000e-04 2.6100e-08 0.0000e+00
+ 2.6240e-08 0.0000e+00 2.6265e-08 6.7000e-04 2.6300e-08 0.0000e+00
+ 2.6440e-08 0.0000e+00 2.6465e-08 6.7000e-04 2.6500e-08 0.0000e+00
+ 2.6640e-08 0.0000e+00 2.6665e-08 6.7000e-04 2.6700e-08 0.0000e+00
+ 2.6840e-08 0.0000e+00 2.6865e-08 6.7000e-04 2.6900e-08 0.0000e+00
+ 2.7040e-08 0.0000e+00 2.7065e-08 6.7000e-04 2.7100e-08 0.0000e+00
+ 2.7240e-08 0.0000e+00 2.7265e-08 6.7000e-04 2.7300e-08 0.0000e+00
+ 2.7440e-08 0.0000e+00 2.7465e-08 6.7000e-04 2.7500e-08 0.0000e+00
+ 2.7640e-08 0.0000e+00 2.7665e-08 6.7000e-04 2.7700e-08 0.0000e+00
+ 2.7840e-08 0.0000e+00 2.7865e-08 6.7000e-04 2.7900e-08 0.0000e+00
+ 2.8040e-08 0.0000e+00 2.8065e-08 6.7000e-04 2.8100e-08 0.0000e+00
+ 2.8240e-08 0.0000e+00 2.8265e-08 6.7000e-04 2.8300e-08 0.0000e+00
+ 2.8440e-08 0.0000e+00 2.8465e-08 6.7000e-04 2.8500e-08 0.0000e+00
+ 2.8640e-08 0.0000e+00 2.8665e-08 6.7000e-04 2.8700e-08 0.0000e+00
+ 2.8840e-08 0.0000e+00 2.8865e-08 6.7000e-04 2.8900e-08 0.0000e+00
+ 2.9040e-08 0.0000e+00 2.9065e-08 6.7000e-04 2.9100e-08 0.0000e+00
+ 2.9240e-08 0.0000e+00 2.9265e-08 6.7000e-04 2.9300e-08 0.0000e+00
+ 2.9440e-08 0.0000e+00 2.9465e-08 6.7000e-04 2.9500e-08 0.0000e+00
+ 2.9640e-08 0.0000e+00 2.9665e-08 6.7000e-04 2.9700e-08 0.0000e+00
+ 2.9840e-08 0.0000e+00 2.9865e-08 6.7000e-04 2.9900e-08 0.0000e+00
+ 3.0040e-08 0.0000e+00 3.0065e-08 6.7000e-04 3.0100e-08 0.0000e+00
+ 3.0240e-08 0.0000e+00 3.0265e-08 6.7000e-04 3.0300e-08 0.0000e+00
+ 3.0440e-08 0.0000e+00 3.0465e-08 6.7000e-04 3.0500e-08 0.0000e+00
+ 3.0640e-08 0.0000e+00 3.0665e-08 6.7000e-04 3.0700e-08 0.0000e+00
+ 3.0840e-08 0.0000e+00 3.0865e-08 6.7000e-04 3.0900e-08 0.0000e+00
+ 3.1040e-08 0.0000e+00 3.1065e-08 6.7000e-04 3.1100e-08 0.0000e+00
+ 3.1240e-08 0.0000e+00 3.1265e-08 6.7000e-04 3.1300e-08 0.0000e+00
+ 3.1440e-08 0.0000e+00 3.1465e-08 6.7000e-04 3.1500e-08 0.0000e+00
+ 3.1640e-08 0.0000e+00 3.1665e-08 6.7000e-04 3.1700e-08 0.0000e+00
+ 3.1840e-08 0.0000e+00 3.1865e-08 6.7000e-04 3.1900e-08 0.0000e+00
+ 3.2040e-08 0.0000e+00 3.2065e-08 6.7000e-04 3.2100e-08 0.0000e+00
+ 3.2240e-08 0.0000e+00 3.2265e-08 6.7000e-04 3.2300e-08 0.0000e+00
+ 3.2440e-08 0.0000e+00 3.2465e-08 6.7000e-04 3.2500e-08 0.0000e+00
+ 3.2640e-08 0.0000e+00 3.2665e-08 6.7000e-04 3.2700e-08 0.0000e+00
+ 3.2840e-08 0.0000e+00 3.2865e-08 6.7000e-04 3.2900e-08 0.0000e+00
+ 3.3040e-08 0.0000e+00 3.3065e-08 6.7000e-04 3.3100e-08 0.0000e+00
+ 3.3240e-08 0.0000e+00 3.3265e-08 6.7000e-04 3.3300e-08 0.0000e+00
+ 3.3440e-08 0.0000e+00 3.3465e-08 6.7000e-04 3.3500e-08 0.0000e+00
+ 3.3640e-08 0.0000e+00 3.3665e-08 6.7000e-04 3.3700e-08 0.0000e+00
+ 3.3840e-08 0.0000e+00 3.3865e-08 6.7000e-04 3.3900e-08 0.0000e+00
+ 3.4040e-08 0.0000e+00 3.4065e-08 6.7000e-04 3.4100e-08 0.0000e+00
+ 3.4240e-08 0.0000e+00 3.4265e-08 6.7000e-04 3.4300e-08 0.0000e+00
+ 3.4440e-08 0.0000e+00 3.4465e-08 6.7000e-04 3.4500e-08 0.0000e+00
+ 3.4640e-08 0.0000e+00 3.4665e-08 6.7000e-04 3.4700e-08 0.0000e+00
+ 3.4840e-08 0.0000e+00 3.4865e-08 6.7000e-04 3.4900e-08 0.0000e+00
+ 3.5040e-08 0.0000e+00 3.5065e-08 6.7000e-04 3.5100e-08 0.0000e+00
+ 3.5240e-08 0.0000e+00 3.5265e-08 6.7000e-04 3.5300e-08 0.0000e+00
+ 3.5440e-08 0.0000e+00 3.5465e-08 6.7000e-04 3.5500e-08 0.0000e+00
+ 3.5640e-08 0.0000e+00 3.5665e-08 6.7000e-04 3.5700e-08 0.0000e+00
+ 3.5840e-08 0.0000e+00 3.5865e-08 6.7000e-04 3.5900e-08 0.0000e+00
+ 3.6040e-08 0.0000e+00 3.6065e-08 6.7000e-04 3.6100e-08 0.0000e+00
+ 3.6240e-08 0.0000e+00 3.6265e-08 6.7000e-04 3.6300e-08 0.0000e+00
+ 3.6440e-08 0.0000e+00 3.6465e-08 6.7000e-04 3.6500e-08 0.0000e+00
+ 3.6640e-08 0.0000e+00 3.6665e-08 6.7000e-04 3.6700e-08 0.0000e+00
+ 3.6840e-08 0.0000e+00 3.6865e-08 6.7000e-04 3.6900e-08 0.0000e+00
+ 3.7040e-08 0.0000e+00 3.7065e-08 6.7000e-04 3.7100e-08 0.0000e+00
+ 3.7240e-08 0.0000e+00 3.7265e-08 6.7000e-04 3.7300e-08 0.0000e+00
+ 3.7440e-08 0.0000e+00 3.7465e-08 6.7000e-04 3.7500e-08 0.0000e+00
+ 3.7640e-08 0.0000e+00 3.7665e-08 6.7000e-04 3.7700e-08 0.0000e+00
+ 3.7840e-08 0.0000e+00 3.7865e-08 6.7000e-04 3.7900e-08 0.0000e+00
+ 3.8040e-08 0.0000e+00 3.8065e-08 6.7000e-04 3.8100e-08 0.0000e+00
+ 3.8240e-08 0.0000e+00 3.8265e-08 6.7000e-04 3.8300e-08 0.0000e+00
+ 3.8440e-08 0.0000e+00 3.8465e-08 6.7000e-04 3.8500e-08 0.0000e+00
+ 3.8640e-08 0.0000e+00 3.8665e-08 6.7000e-04 3.8700e-08 0.0000e+00
+ 3.8840e-08 0.0000e+00 3.8865e-08 6.7000e-04 3.8900e-08 0.0000e+00
+ 3.9040e-08 0.0000e+00 3.9065e-08 6.7000e-04 3.9100e-08 0.0000e+00
+ 3.9240e-08 0.0000e+00 3.9265e-08 6.7000e-04 3.9300e-08 0.0000e+00
+ 3.9440e-08 0.0000e+00 3.9465e-08 6.7000e-04 3.9500e-08 0.0000e+00
+ 3.9640e-08 0.0000e+00 3.9665e-08 6.7000e-04 3.9700e-08 0.0000e+00
+ 3.9840e-08 0.0000e+00 3.9865e-08 6.7000e-04 3.9900e-08 0.0000e+00
+ 4.0040e-08 0.0000e+00 4.0065e-08 6.7000e-04 4.0100e-08 0.0000e+00
+ 4.0240e-08 0.0000e+00 4.0265e-08 6.7000e-04 4.0300e-08 0.0000e+00
+ 4.0440e-08 0.0000e+00 4.0465e-08 6.7000e-04 4.0500e-08 0.0000e+00
+ 4.0640e-08 0.0000e+00 4.0665e-08 6.7000e-04 4.0700e-08 0.0000e+00
+ 4.0840e-08 0.0000e+00 4.0865e-08 6.7000e-04 4.0900e-08 0.0000e+00
+ 4.1040e-08 0.0000e+00 4.1065e-08 6.7000e-04 4.1100e-08 0.0000e+00
+ 4.1240e-08 0.0000e+00 4.1265e-08 6.7000e-04 4.1300e-08 0.0000e+00
+ 4.1440e-08 0.0000e+00 4.1465e-08 6.7000e-04 4.1500e-08 0.0000e+00
+ 4.1640e-08 0.0000e+00 4.1665e-08 6.7000e-04 4.1700e-08 0.0000e+00
+ 4.1840e-08 0.0000e+00 4.1865e-08 6.7000e-04 4.1900e-08 0.0000e+00
+ 4.2040e-08 0.0000e+00 4.2065e-08 6.7000e-04 4.2100e-08 0.0000e+00
+ 4.2240e-08 0.0000e+00 4.2265e-08 6.7000e-04 4.2300e-08 0.0000e+00
+ 4.2440e-08 0.0000e+00 4.2465e-08 6.7000e-04 4.2500e-08 0.0000e+00
+ 4.2640e-08 0.0000e+00 4.2665e-08 6.7000e-04 4.2700e-08 0.0000e+00
+ 4.2840e-08 0.0000e+00 4.2865e-08 6.7000e-04 4.2900e-08 0.0000e+00
+ 4.3040e-08 0.0000e+00 4.3065e-08 6.7000e-04 4.3100e-08 0.0000e+00
+ 4.3240e-08 0.0000e+00 4.3265e-08 6.7000e-04 4.3300e-08 0.0000e+00
+ 4.3440e-08 0.0000e+00 4.3465e-08 6.7000e-04 4.3500e-08 0.0000e+00
+ 4.3640e-08 0.0000e+00 4.3665e-08 6.7000e-04 4.3700e-08 0.0000e+00
+ 4.3840e-08 0.0000e+00 4.3865e-08 6.7000e-04 4.3900e-08 0.0000e+00
+ 4.4040e-08 0.0000e+00 4.4065e-08 6.7000e-04 4.4100e-08 0.0000e+00
+ 4.4240e-08 0.0000e+00 4.4265e-08 6.7000e-04 4.4300e-08 0.0000e+00
+ 4.4440e-08 0.0000e+00 4.4465e-08 6.7000e-04 4.4500e-08 0.0000e+00
+ 4.4640e-08 0.0000e+00 4.4665e-08 6.7000e-04 4.4700e-08 0.0000e+00
+ 4.4840e-08 0.0000e+00 4.4865e-08 6.7000e-04 4.4900e-08 0.0000e+00
+ 4.5040e-08 0.0000e+00 4.5065e-08 6.7000e-04 4.5100e-08 0.0000e+00
+ 4.5240e-08 0.0000e+00 4.5265e-08 6.7000e-04 4.5300e-08 0.0000e+00
+ 4.5440e-08 0.0000e+00 4.5465e-08 6.7000e-04 4.5500e-08 0.0000e+00
+ 4.5640e-08 0.0000e+00 4.5665e-08 6.7000e-04 4.5700e-08 0.0000e+00
+ 4.5840e-08 0.0000e+00 4.5865e-08 6.7000e-04 4.5900e-08 0.0000e+00
+ 4.6040e-08 0.0000e+00 4.6065e-08 6.7000e-04 4.6100e-08 0.0000e+00
+ 4.6240e-08 0.0000e+00 4.6265e-08 6.7000e-04 4.6300e-08 0.0000e+00
+ 4.6440e-08 0.0000e+00 4.6465e-08 6.7000e-04 4.6500e-08 0.0000e+00
+ 4.6640e-08 0.0000e+00 4.6665e-08 6.7000e-04 4.6700e-08 0.0000e+00
+ 4.6840e-08 0.0000e+00 4.6865e-08 6.7000e-04 4.6900e-08 0.0000e+00
+ 4.7040e-08 0.0000e+00 4.7065e-08 6.7000e-04 4.7100e-08 0.0000e+00
+ 4.7240e-08 0.0000e+00 4.7265e-08 6.7000e-04 4.7300e-08 0.0000e+00
+ 4.7440e-08 0.0000e+00 4.7465e-08 6.7000e-04 4.7500e-08 0.0000e+00
+ 4.7640e-08 0.0000e+00 4.7665e-08 6.7000e-04 4.7700e-08 0.0000e+00
+ 4.7840e-08 0.0000e+00 4.7865e-08 6.7000e-04 4.7900e-08 0.0000e+00
+ 4.8040e-08 0.0000e+00 4.8065e-08 6.7000e-04 4.8100e-08 0.0000e+00
+ 4.8240e-08 0.0000e+00 4.8265e-08 6.7000e-04 4.8300e-08 0.0000e+00
+ 4.8440e-08 0.0000e+00 4.8465e-08 6.7000e-04 4.8500e-08 0.0000e+00
+ 4.8640e-08 0.0000e+00 4.8665e-08 6.7000e-04 4.8700e-08 0.0000e+00
+ 4.8840e-08 0.0000e+00 4.8865e-08 6.7000e-04 4.8900e-08 0.0000e+00
+ 4.9040e-08 0.0000e+00 4.9065e-08 6.7000e-04 4.9100e-08 0.0000e+00
+ 4.9240e-08 0.0000e+00 4.9265e-08 6.7000e-04 4.9300e-08 0.0000e+00
+ 4.9440e-08 0.0000e+00 4.9465e-08 6.7000e-04 4.9500e-08 0.0000e+00
+ 4.9640e-08 0.0000e+00 4.9665e-08 6.7000e-04 4.9700e-08 0.0000e+00
+ 4.9840e-08 0.0000e+00 4.9865e-08 6.7000e-04 4.9900e-08 0.0000e+00
+ 5.0040e-08 0.0000e+00 5.0065e-08 6.7000e-04 5.0100e-08 0.0000e+00
+ 5.0240e-08 0.0000e+00 5.0265e-08 6.7000e-04 5.0300e-08 0.0000e+00
+ 5.0440e-08 0.0000e+00 5.0465e-08 6.7000e-04 5.0500e-08 0.0000e+00
+ 5.0640e-08 0.0000e+00 5.0665e-08 6.7000e-04 5.0700e-08 0.0000e+00
+ 5.0840e-08 0.0000e+00 5.0865e-08 6.7000e-04 5.0900e-08 0.0000e+00
+ 5.1040e-08 0.0000e+00 5.1065e-08 6.7000e-04 5.1100e-08 0.0000e+00
+ 5.1240e-08 0.0000e+00 5.1265e-08 6.7000e-04 5.1300e-08 0.0000e+00
+ 5.1440e-08 0.0000e+00 5.1465e-08 6.7000e-04 5.1500e-08 0.0000e+00
+ 5.1640e-08 0.0000e+00 5.1665e-08 6.7000e-04 5.1700e-08 0.0000e+00
+ 5.1840e-08 0.0000e+00 5.1865e-08 6.7000e-04 5.1900e-08 0.0000e+00
+ 5.2040e-08 0.0000e+00 5.2065e-08 6.7000e-04 5.2100e-08 0.0000e+00
+ 5.2240e-08 0.0000e+00 5.2265e-08 6.7000e-04 5.2300e-08 0.0000e+00
+ 5.2440e-08 0.0000e+00 5.2465e-08 6.7000e-04 5.2500e-08 0.0000e+00
+ 5.2640e-08 0.0000e+00 5.2665e-08 6.7000e-04 5.2700e-08 0.0000e+00
+ 5.2840e-08 0.0000e+00 5.2865e-08 6.7000e-04 5.2900e-08 0.0000e+00
+ 5.3040e-08 0.0000e+00 5.3065e-08 6.7000e-04 5.3100e-08 0.0000e+00
+ 5.3240e-08 0.0000e+00 5.3265e-08 6.7000e-04 5.3300e-08 0.0000e+00
+ 5.3440e-08 0.0000e+00 5.3465e-08 6.7000e-04 5.3500e-08 0.0000e+00
+ 5.3640e-08 0.0000e+00 5.3665e-08 6.7000e-04 5.3700e-08 0.0000e+00
+ 5.3840e-08 0.0000e+00 5.3865e-08 6.7000e-04 5.3900e-08 0.0000e+00
+ 5.4040e-08 0.0000e+00 5.4065e-08 6.7000e-04 5.4100e-08 0.0000e+00
+ 5.4240e-08 0.0000e+00 5.4265e-08 6.7000e-04 5.4300e-08 0.0000e+00
+ 5.4440e-08 0.0000e+00 5.4465e-08 6.7000e-04 5.4500e-08 0.0000e+00
+ 5.4640e-08 0.0000e+00 5.4665e-08 6.7000e-04 5.4700e-08 0.0000e+00
+ 5.4840e-08 0.0000e+00 5.4865e-08 6.7000e-04 5.4900e-08 0.0000e+00
+ 5.5040e-08 0.0000e+00 5.5065e-08 6.7000e-04 5.5100e-08 0.0000e+00
+ 5.5240e-08 0.0000e+00 5.5265e-08 6.7000e-04 5.5300e-08 0.0000e+00
+ 5.5440e-08 0.0000e+00 5.5465e-08 6.7000e-04 5.5500e-08 0.0000e+00
+ 5.5640e-08 0.0000e+00 5.5665e-08 6.7000e-04 5.5700e-08 0.0000e+00
+ 5.5840e-08 0.0000e+00 5.5865e-08 6.7000e-04 5.5900e-08 0.0000e+00
+ 5.6040e-08 0.0000e+00 5.6065e-08 6.7000e-04 5.6100e-08 0.0000e+00
+ 5.6240e-08 0.0000e+00 5.6265e-08 6.7000e-04 5.6300e-08 0.0000e+00
+ 5.6440e-08 0.0000e+00 5.6465e-08 6.7000e-04 5.6500e-08 0.0000e+00
+ 5.6640e-08 0.0000e+00 5.6665e-08 6.7000e-04 5.6700e-08 0.0000e+00
+ 5.6840e-08 0.0000e+00 5.6865e-08 6.7000e-04 5.6900e-08 0.0000e+00
+ 5.7040e-08 0.0000e+00 5.7065e-08 6.7000e-04 5.7100e-08 0.0000e+00
+ 5.7240e-08 0.0000e+00 5.7265e-08 6.7000e-04 5.7300e-08 0.0000e+00
+ 5.7440e-08 0.0000e+00 5.7465e-08 6.7000e-04 5.7500e-08 0.0000e+00
+ 5.7640e-08 0.0000e+00 5.7665e-08 6.7000e-04 5.7700e-08 0.0000e+00
+ 5.7840e-08 0.0000e+00 5.7865e-08 6.7000e-04 5.7900e-08 0.0000e+00
+ 5.8040e-08 0.0000e+00 5.8065e-08 6.7000e-04 5.8100e-08 0.0000e+00
+ 5.8240e-08 0.0000e+00 5.8265e-08 6.7000e-04 5.8300e-08 0.0000e+00
+ 5.8440e-08 0.0000e+00 5.8465e-08 6.7000e-04 5.8500e-08 0.0000e+00
+ 5.8640e-08 0.0000e+00 5.8665e-08 6.7000e-04 5.8700e-08 0.0000e+00
+ 5.8840e-08 0.0000e+00 5.8865e-08 6.7000e-04 5.8900e-08 0.0000e+00
+ 5.9040e-08 0.0000e+00 5.9065e-08 6.7000e-04 5.9100e-08 0.0000e+00
+ 5.9240e-08 0.0000e+00 5.9265e-08 6.7000e-04 5.9300e-08 0.0000e+00
+ 5.9440e-08 0.0000e+00 5.9465e-08 6.7000e-04 5.9500e-08 0.0000e+00
+ 5.9640e-08 0.0000e+00 5.9665e-08 6.7000e-04 5.9700e-08 0.0000e+00
+ 5.9840e-08 0.0000e+00 5.9865e-08 6.7000e-04 5.9900e-08 0.0000e+00
+ 6.0040e-08 0.0000e+00 6.0065e-08 6.7000e-04 6.0100e-08 0.0000e+00
+ 6.0240e-08 0.0000e+00 6.0265e-08 6.7000e-04 6.0300e-08 0.0000e+00
+ 6.0440e-08 0.0000e+00 6.0465e-08 6.7000e-04 6.0500e-08 0.0000e+00)

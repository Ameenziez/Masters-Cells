
#works well!
#got the data to propagate
.include LSmitll_DCSFQ_PTLTX_v1p5.cir
.include LSmitll_bufft_v1p5.cir
.include LSmitll_PTLRX_SFQDC_v1p5.cir
.include LSmitll_SPLITT_v1p5.cir
.INCLUDE LSMITLL_JTLT_V1P5.CIR
.INCLUDE LSMITLL_MERGET_V1P5.CIR
.include storeedit.cir
.INCLUDE COMPONENTSEDIT.CIR
.INCLUDE COMP3.CIR
.INCLUDE COMP4.CIR
.INCLUDE COMP5.CIR
.include conv.cir
.INCLUDE synapsenext2.CIR
.INCLUDE DCPULSER.CIR
.INCLUDE MULTISPLIT.CIR
.include transmit.cir
.INCLUDE DELAY7.CIR
.INCLUDE AND.CIR
.INCLUDE AND3.CIR
.INCLUDE OR3.CIR
.include PERCEPTRON.CIR
.include CONVINTERFACE.cir
.INCLUDE COMP6.CIR


# TRY SHIFTING CLK OF OUTPUT BACK A BIT...
#.tran 1ps 45000PS 0ps 1p
.tran 1ps 15000PS 0ps 1p
#MLP:
#D=Oi.T + Oi.!Oj + T.!Oj 

#setup circuitry
#VAC1   A1   0   SIN(0 723mV 10GHz 200Ps 0)
VAC1   A1   0   SIN(0 723mV 10GHz 400Ps 0)
RAC1   A1   A2   1000
LAC1   A2   A3   0.1p
#VAC2   B1   0   SIN(0 723mV 10GHz 175.0ps 0)
VAC2   B1   0   SIN(0 723mV 10GHz 375.0ps 0)
RAC2   B1   B2   1000
LAC2   B2   B3   0.1p
VDC    DC1   0   pwl(0 0 20p 1023mV)
RDC    DC1   DC2   1000
LDC    DC2   DC3  0.1p
VDCconv    DCc1   0   PWL(0ps 0mV 20ps 1023mV 60000p 1023mV 60000p 0)
#was 640
RDCconv    DCc1   DCc2  640
LDCconv    DCc2   DCc3   0.1p


LTARGET1 TARGET0 TARGET1 1p

#SPLIT INPUTS BETWEEN 2 NEURONS
LINPUT1 IN1 INPUT11 1P
LINPUT2 IN2 INPUT12 1P
LINPUTBIAS11 INB11 INPUTB 1P

#3,-1,1 works
.param flx1=3
.param flx2=-1
.param flxb=1
#.param flx1=-2
#.param flx2=0
#.param flxb=1
#.param flx1=-1
#.param flx2=1
#.param flxb=2

IINITAL11 0 INITIAL11 PWL( 0 0 20P -22.3U*flx1 3000p -22.3U*flx1 3001p 0 )
IINITAL12 0 INITIAL12 PWL( 0 0 20P -22.3U*flx2 3000p -22.3U*flx2 3001p 0)
IINITALB11 0 INITIALB11 PWL( 0 0 20P -22.3u*flxb 3000p -22.3U*flxb 3001p 0)

#IINITAL11 0 INITIAL11 PWL( 0 0 20P -22.3U*flx1  )
#IINITAL12 0 INITIAL12 PWL( 0 0 20P -22.3U*flx2 )
#IINITALB11 0 INITIALB11 PWL( 0 0 20P -22.3u*flxb )




##FINAL ACTIVATION - this works 
ITHRESH11 0 THRESH11 PWL(0 0 20p 10U)

#buffers for input and target

XNEURON 3NEURON2 INPUT11 INPUT12 INPUTB TARGET1  THRESH11 A3 0 B3 0 DC3 0 DCC3 0 INITIAL11 INITIAL12 INITIALB11
          #x3NEURON2 INPUT1 INPUT2 INPUTBIAS TARGET DOUTFINAL1 DOUTFINAL2 THRESH XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT DCCIN DCCOUT OUTPUT OUTPUTAXON











.PRINT DEVII IIN1
.PRINT DEVII IIN2
#.PRINT DEVII IINBIAS1
.PRINT DEVII ITARGET
.print phase lq.XACT.XNEURON

#.print phase LQ.X11.XNEURON
#.print phase LQ.X12.XNEURON
#.print phase lQ.XB11.XNEURON

#.print phase lstore1.X11.XNEURON
#.print phase lstore1.X12.XNEURON
#.print phase lstore1.XB11.XNEURON



#.print phase l1_q.xdecr.XPERCEPTRON11.XNEURON1
#.print phase l2_q.xdecr.XPERCEPTRON11.XNEURON1
#.print phase l4_q.xdecr.XPERCEPTRON11.XNEURON1
#.print phase l5_q.xdecr.XPERCEPTRON11.XNEURON1
#.print phase l5_q.xDEcr.XPERCEPTRON11.XNEURON1


#.print phase lq.xinput.XPERCEPTRONb11.XNEURON1
#.print phase lq.XTARGET.XPERCEPTRONb11.XNEURON1
#.print phase l1_q.xincr.XPERCEPTRONB11.XNEURON1
#.print phase l2_q.xincr.XPERCEPTRONB11.XNEURON1
#.print phase l4_q.xincr.XPERCEPTRONB11.XNEURON1
#.print phase l5_q.xincr.XPERCEPTRONB11.XNEURON1

#.print phase l1_q.xDEcr.XPERCEPTRONb11.XNEURON1
#.print phase l2_q.xDEcr.XPERCEPTRONb11.XNEURON1
#.print phase l4_q.xDEcr.XPERCEPTRONb11.XNEURON1
#.print phase l5_q.xDEcr.XPERCEPTRONb11.XNEURON1










.SUBCKT 3NEURON2 INPUT1 INPUT2 INPUTBIAS TARGET THRESH XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT DCCIN DCCOUT INITIAL11 INITIAL12 INITIALB11

#INPUTS
LSYN11 INPUT1 SYN11 1p  
LSYN12 INPUT2 SYN12 1p  
LSYNB11 INPUTBIAS SYNB11 1p  
LTARGET1 TARGET TARGET1 1p
LTARGET2 TARGET1 0 1p

#COUPLINGS
KSYN11 LSYN11 LSYNADJUST11 -0.05
KSYN12 LSYN12 LSYNADJUST12 -0.05
KSYNB11 LSYNB11 LSYNADJUSTB11 -0.05
KT1 LTARGET1 LADJUSTTARGET1 -0.05
LSYNADJUST11 0 ADJUST11 5P 
LSYNADJUST12 0 ADJUST12 5P 
LSYNADJUSTB11 0 ADJUSTB11 5P 
LADJUSTTARGET1 0 ADJUSTTARGET1 5P


#SYNAPSE 1
XSTORE11 BISTORE SFQOUTPLUS11 SFQOUTMINUS11 WEIGHTL11 WEIGHTR11
X11 SYNAPSEfastest SYN11 DOUT12 DOUT11 WEIGHTL11 WEIGHTR11 INITIAL11


#SYNAPSE 2
XSTORE12 BISTORE SFQOUTPLUS12 SFQOUTMINUS12 WEIGHTL12 WEIGHTR12
X12 SYNAPSEfastest SYN12 DOUT13 DOUT12 WEIGHTL12 WEIGHTR12 INITIAL12

#SYNAPSE BIAS
XSTOREB11 BISTORE SFQOUTPLUSB11 SFQOUTMINUSB11 WEIGHTLB11 WEIGHTRB11
XB11 SYNAPSEfastest SYNB11 0 DOUT13 WEIGHTLB11 WEIGHTRB11 INITIALB11

#ACTIVATION
XACT COMP6 XIN1 DOUT11 A4 DCIN DC4 DOUTL11 0  0 DOUTR12   DOUTL13 0 0 DOUTR14   DOUTL15 0 0 DOUTR16   THRESH


#DELAYS
XTARGETDELAY bfrsplit3 A4 ADJUSTTARGET1 A5 DC4 DC5 0 TARGETDELAYED1 0 TARGETDELAYED2 0 TARGETDELAYED3
XINPUT1DELAY BFR A5 ADJUST11 A6 DC5 DC6 0 INPUT1DELAYED
XINPUT2DELAY BFR A6 ADJUST12 A7 DC6 DC7 0 INPUT2DELAYED
XINPUTB1DELAY BFR A7 ADJUSTB11 A14 DC7 DC14 0 INPUTB1DELAYED



#XPERCEPTRON11 PERCEPTRON  B13 XIN2  A14 A15  INPUT1DELAYED DOUTL11 DOUTR12  TARGETDELAYED1 DC15 DC14 INCR11 DECR11
#XPERCEPTRON12 PERCEPTRON  B14 B13  A15 A16  INPUT2DELAYED DOUTL13 DOUTR14 TARGETDELAYED2 DC16 DC15 INCR12 DECR12
#XPERCEPTRONB11 PERCEPTRON  XOUT2 B14  A16 A17  INPUTB1DELAYED DOUTL15 DOUTR16 TARGETDELAYED3 DCOUT DC16 INCRB11 DECRB11



#XCONV11 CONV A17 A18 DCC5 DCCIN INCR11 DECR11 SFQOUTPLUS11 SFQOUTMINUS11
#XCONV12 CONV A18 A19 DCC6 DCC5 INCR12 DECR12 SFQOUTPLUS12 SFQOUTMINUS12
#XCONVB11 CONV A19 XOUT1 DCCOUT DCC6 INCRB11 DECRB11 SFQOUTPLUSB11 SFQOUTMINUSB11

######TINKERED FROM HERE####
XPERCEPTRON11 PERCEPTRON  B13 XIN2  A14 A15  INPUT1DELAYED  DOUTR12 DOUTL11 TARGETDELAYED1 DC15 DC14 INCR11 DECR11
XPERCEPTRON12 PERCEPTRON  B14 B13  A15 A16  INPUT2DELAYED  DOUTR14 DOUTL13 TARGETDELAYED2 DC16 DC15 INCR12 DECR12
XPERCEPTRONB11 PERCEPTRON  XOUT2 B14  A16 A17  INPUTB1DELAYED  DOUTR16 DOUTL15 TARGETDELAYED3 DCOUT DC16 INCRB11 DECRB11
#SWITCHED INCR AND DECR BECAUSE FOR SOME REASON IT GOT SWITCHED...


XCONV11 CONV A17 A18 DCC5 DCCIN DECR11 INCR11  SFQOUTPLUS11 SFQOUTMINUS11
XCONV12 CONV A18 A19 DCC6 DCC5 DECR12 INCR12  SFQOUTPLUS12 SFQOUTMINUS12
XCONVB11 CONV A19 XOUT1 DCCOUT DCC6  DECRB11 INCRB11 SFQOUTPLUSB11 SFQOUTMINUSB11

.ENDS 3NEURON2











***    INPUTS  ***
IIN1 0 IN1 PWL(0 0 20P 0 7.5000e-10 0.0000e+00 7.5500e-10 1.0000e-03 8.0500e-10 1.0000e-03
+ 8.1000e-10 0.0000e+00 1.1500e-09 0.0000e+00 1.1550e-09 1.0000e-03
+ 1.2050e-09 1.0000e-03 1.2100e-09 0.0000e+00 1.5500e-09 0.0000e+00
+ 1.5550e-09 1.0000e-03 1.6050e-09 1.0000e-03 1.6100e-09 0.0000e+00
+ 1.9500e-09 0.0000e+00 1.9550e-09 1.0000e-03 2.0050e-09 1.0000e-03
+ 2.0100e-09 0.0000e+00 2.3500e-09 0.0000e+00 2.3550e-09 1.0000e-03
+ 2.4050e-09 1.0000e-03 2.4100e-09 0.0000e+00 2.7500e-09 0.0000e+00
+ 2.7550e-09 1.0000e-03 2.8050e-09 1.0000e-03 2.8100e-09 0.0000e+00
+ 3.1500e-09 0.0000e+00 3.1550e-09 1.0000e-03 3.2050e-09 1.0000e-03
+ 3.2100e-09 0.0000e+00 3.5500e-09 0.0000e+00 3.5550e-09 1.0000e-03
+ 3.6050e-09 1.0000e-03 3.6100e-09 0.0000e+00 3.9500e-09 0.0000e+00
+ 3.9550e-09 1.0000e-03 4.0050e-09 1.0000e-03 4.0100e-09 0.0000e+00
+ 4.3500e-09 0.0000e+00 4.3550e-09 1.0000e-03 4.4050e-09 1.0000e-03
+ 4.4100e-09 0.0000e+00 4.7500e-09 0.0000e+00 4.7550e-09 1.0000e-03
+ 4.8050e-09 1.0000e-03 4.8100e-09 0.0000e+00 5.1500e-09 0.0000e+00
+ 5.1550e-09 1.0000e-03 5.2050e-09 1.0000e-03 5.2100e-09 0.0000e+00
+ 5.5500e-09 0.0000e+00 5.5550e-09 1.0000e-03 5.6050e-09 1.0000e-03
+ 5.6100e-09 0.0000e+00 5.9500e-09 0.0000e+00 5.9550e-09 1.0000e-03
+ 6.0050e-09 1.0000e-03 6.0100e-09 0.0000e+00 6.3500e-09 0.0000e+00
+ 6.3550e-09 1.0000e-03 6.4050e-09 1.0000e-03 6.4100e-09 0.0000e+00
+ 6.7500e-09 0.0000e+00 6.7550e-09 1.0000e-03 6.8050e-09 1.0000e-03
+ 6.8100e-09 0.0000e+00 7.1500e-09 0.0000e+00 7.1550e-09 1.0000e-03
+ 7.2050e-09 1.0000e-03 7.2100e-09 0.0000e+00 7.5500e-09 0.0000e+00
+ 7.5550e-09 1.0000e-03 7.6050e-09 1.0000e-03 7.6100e-09 0.0000e+00
+ 7.9500e-09 0.0000e+00 7.9550e-09 1.0000e-03 8.0050e-09 1.0000e-03
+ 8.0100e-09 0.0000e+00 8.3500e-09 0.0000e+00 8.3550e-09 1.0000e-03
+ 8.4050e-09 1.0000e-03 8.4100e-09 0.0000e+00 8.7500e-09 0.0000e+00
+ 8.7550e-09 1.0000e-03 8.8050e-09 1.0000e-03 8.8100e-09 0.0000e+00
+ 9.1500e-09 0.0000e+00 9.1550e-09 1.0000e-03 9.2050e-09 1.0000e-03
+ 9.2100e-09 0.0000e+00 9.5500e-09 0.0000e+00 9.5550e-09 1.0000e-03
+ 9.6050e-09 1.0000e-03 9.6100e-09 0.0000e+00 9.9500e-09 0.0000e+00
+ 9.9550e-09 1.0000e-03 1.0005e-08 1.0000e-03 1.0010e-08 0.0000e+00
+ 1.0350e-08 0.0000e+00 1.0355e-08 1.0000e-03 1.0405e-08 1.0000e-03
+ 1.0410e-08 0.0000e+00 1.0750e-08 0.0000e+00 1.0755e-08 1.0000e-03
+ 1.0805e-08 1.0000e-03 1.0810e-08 0.0000e+00 1.1150e-08 0.0000e+00
+ 1.1155e-08 1.0000e-03 1.1205e-08 1.0000e-03 1.1210e-08 0.0000e+00
+ 1.1550e-08 0.0000e+00 1.1555e-08 1.0000e-03 1.1605e-08 1.0000e-03
+ 1.1610e-08 0.0000e+00 1.1950e-08 0.0000e+00 1.1955e-08 1.0000e-03
+ 1.2005e-08 1.0000e-03 1.2010e-08 0.0000e+00 1.2350e-08 0.0000e+00
+ 1.2355e-08 1.0000e-03 1.2405e-08 1.0000e-03 1.2410e-08 0.0000e+00
+ 1.2750e-08 0.0000e+00 1.2755e-08 1.0000e-03 1.2805e-08 1.0000e-03
+ 1.2810e-08 0.0000e+00 1.3150e-08 0.0000e+00 1.3155e-08 1.0000e-03
+ 1.3205e-08 1.0000e-03 1.3210e-08 0.0000e+00 1.3550e-08 0.0000e+00
+ 1.3555e-08 1.0000e-03 1.3605e-08 1.0000e-03 1.3610e-08 0.0000e+00
+ 1.3950e-08 0.0000e+00 1.3955e-08 1.0000e-03 1.4005e-08 1.0000e-03
+ 1.4010e-08 0.0000e+00 1.4350e-08 0.0000e+00 1.4355e-08 1.0000e-03
+ 1.4405e-08 1.0000e-03 1.4410e-08 0.0000e+00 1.4750e-08 0.0000e+00
+ 1.4755e-08 1.0000e-03 1.4805e-08 1.0000e-03 1.4810e-08 0.0000e+00
+ 1.5150e-08 0.0000e+00 1.5155e-08 1.0000e-03 1.5205e-08 1.0000e-03
+ 1.5210e-08 0.0000e+00 1.5550e-08 0.0000e+00 1.5555e-08 1.0000e-03
+ 1.5605e-08 1.0000e-03 1.5610e-08 0.0000e+00 1.5950e-08 0.0000e+00
+ 1.5955e-08 1.0000e-03 1.6005e-08 1.0000e-03 1.6010e-08 0.0000e+00
+ 1.6350e-08 0.0000e+00 1.6355e-08 1.0000e-03 1.6405e-08 1.0000e-03
+ 1.6410e-08 0.0000e+00 1.6750e-08 0.0000e+00 1.6755e-08 1.0000e-03
+ 1.6805e-08 1.0000e-03 1.6810e-08 0.0000e+00 1.7150e-08 0.0000e+00
+ 1.7155e-08 1.0000e-03 1.7205e-08 1.0000e-03 1.7210e-08 0.0000e+00
+ 1.7550e-08 0.0000e+00 1.7555e-08 1.0000e-03 1.7605e-08 1.0000e-03
+ 1.7610e-08 0.0000e+00 1.7950e-08 0.0000e+00 1.7955e-08 1.0000e-03
+ 1.8005e-08 1.0000e-03 1.8010e-08 0.0000e+00 1.8350e-08 0.0000e+00
+ 1.8355e-08 1.0000e-03 1.8405e-08 1.0000e-03 1.8410e-08 0.0000e+00
+ 1.8750e-08 0.0000e+00 1.8755e-08 1.0000e-03 1.8805e-08 1.0000e-03
+ 1.8810e-08 0.0000e+00 1.9150e-08 0.0000e+00 1.9155e-08 1.0000e-03
+ 1.9205e-08 1.0000e-03 1.9210e-08 0.0000e+00 1.9550e-08 0.0000e+00
+ 1.9555e-08 1.0000e-03 1.9605e-08 1.0000e-03 1.9610e-08 0.0000e+00
+ 1.9950e-08 0.0000e+00 1.9955e-08 1.0000e-03 2.0005e-08 1.0000e-03
+ 2.0010e-08 0.0000e+00 2.0350e-08 0.0000e+00 2.0355e-08 1.0000e-03
+ 2.0405e-08 1.0000e-03 2.0410e-08 0.0000e+00 2.0750e-08 0.0000e+00
+ 2.0755e-08 1.0000e-03 2.0805e-08 1.0000e-03 2.0810e-08 0.0000e+00
+ 2.1150e-08 0.0000e+00 2.1155e-08 1.0000e-03 2.1205e-08 1.0000e-03
+ 2.1210e-08 0.0000e+00 2.1550e-08 0.0000e+00 2.1555e-08 1.0000e-03
+ 2.1605e-08 1.0000e-03 2.1610e-08 0.0000e+00 2.1950e-08 0.0000e+00
+ 2.1955e-08 1.0000e-03 2.2005e-08 1.0000e-03 2.2010e-08 0.0000e+00
+ 2.2350e-08 0.0000e+00 2.2355e-08 1.0000e-03 2.2405e-08 1.0000e-03
+ 2.2410e-08 0.0000e+00 2.2750e-08 0.0000e+00 2.2755e-08 1.0000e-03
+ 2.2805e-08 1.0000e-03 2.2810e-08 0.0000e+00 2.3150e-08 0.0000e+00
+ 2.3155e-08 1.0000e-03 2.3205e-08 1.0000e-03 2.3210e-08 0.0000e+00
+ 2.3550e-08 0.0000e+00 2.3555e-08 1.0000e-03 2.3605e-08 1.0000e-03
+ 2.3610e-08 0.0000e+00 2.3950e-08 0.0000e+00 2.3955e-08 1.0000e-03
+ 2.4005e-08 1.0000e-03 2.4010e-08 0.0000e+00 2.4350e-08 0.0000e+00
+ 2.4355e-08 1.0000e-03 2.4405e-08 1.0000e-03 2.4410e-08 0.0000e+00
+ 2.4750e-08 0.0000e+00 2.4755e-08 1.0000e-03 2.4805e-08 1.0000e-03
+ 2.4810e-08 0.0000e+00 2.5150e-08 0.0000e+00 2.5155e-08 1.0000e-03
+ 2.5205e-08 1.0000e-03 2.5210e-08 0.0000e+00 2.5550e-08 0.0000e+00
+ 2.5555e-08 1.0000e-03 2.5605e-08 1.0000e-03 2.5610e-08 0.0000e+00
+ 2.5950e-08 0.0000e+00 2.5955e-08 1.0000e-03 2.6005e-08 1.0000e-03
+ 2.6010e-08 0.0000e+00 2.6350e-08 0.0000e+00 2.6355e-08 1.0000e-03
+ 2.6405e-08 1.0000e-03 2.6410e-08 0.0000e+00 2.6750e-08 0.0000e+00
+ 2.6755e-08 1.0000e-03 2.6805e-08 1.0000e-03 2.6810e-08 0.0000e+00
+ 2.7150e-08 0.0000e+00 2.7155e-08 1.0000e-03 2.7205e-08 1.0000e-03
+ 2.7210e-08 0.0000e+00 2.7550e-08 0.0000e+00 2.7555e-08 1.0000e-03
+ 2.7605e-08 1.0000e-03 2.7610e-08 0.0000e+00 2.7950e-08 0.0000e+00
+ 2.7955e-08 1.0000e-03 2.8005e-08 1.0000e-03 2.8010e-08 0.0000e+00
+ 2.8350e-08 0.0000e+00 2.8355e-08 1.0000e-03 2.8405e-08 1.0000e-03
+ 2.8410e-08 0.0000e+00 2.8750e-08 0.0000e+00 2.8755e-08 1.0000e-03
+ 2.8805e-08 1.0000e-03 2.8810e-08 0.0000e+00 2.9150e-08 0.0000e+00
+ 2.9155e-08 1.0000e-03 2.9205e-08 1.0000e-03 2.9210e-08 0.0000e+00
+ 2.9550e-08 0.0000e+00 2.9555e-08 1.0000e-03 2.9605e-08 1.0000e-03
+ 2.9610e-08 0.0000e+00 2.9950e-08 0.0000e+00 2.9955e-08 1.0000e-03
+ 3.0005e-08 1.0000e-03 3.0010e-08 0.0000e+00 3.0350e-08 0.0000e+00
+ 3.0355e-08 1.0000e-03 3.0405e-08 1.0000e-03 3.0410e-08 0.0000e+00
+ 3.0750e-08 0.0000e+00 3.0755e-08 1.0000e-03 3.0805e-08 1.0000e-03
+ 3.0810e-08 0.0000e+00 3.1150e-08 0.0000e+00 3.1155e-08 1.0000e-03
+ 3.1205e-08 1.0000e-03 3.1210e-08 0.0000e+00 3.1550e-08 0.0000e+00
+ 3.1555e-08 1.0000e-03 3.1605e-08 1.0000e-03 3.1610e-08 0.0000e+00
+ 3.1950e-08 0.0000e+00 3.1955e-08 1.0000e-03 3.2005e-08 1.0000e-03
+ 3.2010e-08 0.0000e+00 3.2350e-08 0.0000e+00 3.2355e-08 1.0000e-03
+ 3.2405e-08 1.0000e-03 3.2410e-08 0.0000e+00)
IIN2 0 IN2 PWL(0 0 20P 0 9.5000e-10 0.0000e+00 9.5500e-10 1.0000e-03 1.0050e-09 1.0000e-03
+ 1.0100e-09 0.0000e+00 1.1500e-09 0.0000e+00 1.1550e-09 1.0000e-03
+ 1.2050e-09 1.0000e-03 1.2100e-09 0.0000e+00 1.7500e-09 0.0000e+00
+ 1.7550e-09 1.0000e-03 1.8050e-09 1.0000e-03 1.8100e-09 0.0000e+00
+ 1.9500e-09 0.0000e+00 1.9550e-09 1.0000e-03 2.0050e-09 1.0000e-03
+ 2.0100e-09 0.0000e+00 2.5500e-09 0.0000e+00 2.5550e-09 1.0000e-03
+ 2.6050e-09 1.0000e-03 2.6100e-09 0.0000e+00 2.7500e-09 0.0000e+00
+ 2.7550e-09 1.0000e-03 2.8050e-09 1.0000e-03 2.8100e-09 0.0000e+00
+ 3.3500e-09 0.0000e+00 3.3550e-09 1.0000e-03 3.4050e-09 1.0000e-03
+ 3.4100e-09 0.0000e+00 3.5500e-09 0.0000e+00 3.5550e-09 1.0000e-03
+ 3.6050e-09 1.0000e-03 3.6100e-09 0.0000e+00 4.1500e-09 0.0000e+00
+ 4.1550e-09 1.0000e-03 4.2050e-09 1.0000e-03 4.2100e-09 0.0000e+00
+ 4.3500e-09 0.0000e+00 4.3550e-09 1.0000e-03 4.4050e-09 1.0000e-03
+ 4.4100e-09 0.0000e+00 4.9500e-09 0.0000e+00 4.9550e-09 1.0000e-03
+ 5.0050e-09 1.0000e-03 5.0100e-09 0.0000e+00 5.1500e-09 0.0000e+00
+ 5.1550e-09 1.0000e-03 5.2050e-09 1.0000e-03 5.2100e-09 0.0000e+00
+ 5.7500e-09 0.0000e+00 5.7550e-09 1.0000e-03 5.8050e-09 1.0000e-03
+ 5.8100e-09 0.0000e+00 5.9500e-09 0.0000e+00 5.9550e-09 1.0000e-03
+ 6.0050e-09 1.0000e-03 6.0100e-09 0.0000e+00 6.5500e-09 0.0000e+00
+ 6.5550e-09 1.0000e-03 6.6050e-09 1.0000e-03 6.6100e-09 0.0000e+00
+ 6.7500e-09 0.0000e+00 6.7550e-09 1.0000e-03 6.8050e-09 1.0000e-03
+ 6.8100e-09 0.0000e+00 7.3500e-09 0.0000e+00 7.3550e-09 1.0000e-03
+ 7.4050e-09 1.0000e-03 7.4100e-09 0.0000e+00 7.5500e-09 0.0000e+00
+ 7.5550e-09 1.0000e-03 7.6050e-09 1.0000e-03 7.6100e-09 0.0000e+00
+ 8.1500e-09 0.0000e+00 8.1550e-09 1.0000e-03 8.2050e-09 1.0000e-03
+ 8.2100e-09 0.0000e+00 8.3500e-09 0.0000e+00 8.3550e-09 1.0000e-03
+ 8.4050e-09 1.0000e-03 8.4100e-09 0.0000e+00 8.9500e-09 0.0000e+00
+ 8.9550e-09 1.0000e-03 9.0050e-09 1.0000e-03 9.0100e-09 0.0000e+00
+ 9.1500e-09 0.0000e+00 9.1550e-09 1.0000e-03 9.2050e-09 1.0000e-03
+ 9.2100e-09 0.0000e+00 9.7500e-09 0.0000e+00 9.7550e-09 1.0000e-03
+ 9.8050e-09 1.0000e-03 9.8100e-09 0.0000e+00 9.9500e-09 0.0000e+00
+ 9.9550e-09 1.0000e-03 1.0005e-08 1.0000e-03 1.0010e-08 0.0000e+00
+ 1.0550e-08 0.0000e+00 1.0555e-08 1.0000e-03 1.0605e-08 1.0000e-03
+ 1.0610e-08 0.0000e+00 1.0750e-08 0.0000e+00 1.0755e-08 1.0000e-03
+ 1.0805e-08 1.0000e-03 1.0810e-08 0.0000e+00 1.1350e-08 0.0000e+00
+ 1.1355e-08 1.0000e-03 1.1405e-08 1.0000e-03 1.1410e-08 0.0000e+00
+ 1.1550e-08 0.0000e+00 1.1555e-08 1.0000e-03 1.1605e-08 1.0000e-03
+ 1.1610e-08 0.0000e+00 1.2150e-08 0.0000e+00 1.2155e-08 1.0000e-03
+ 1.2205e-08 1.0000e-03 1.2210e-08 0.0000e+00 1.2350e-08 0.0000e+00
+ 1.2355e-08 1.0000e-03 1.2405e-08 1.0000e-03 1.2410e-08 0.0000e+00
+ 1.2950e-08 0.0000e+00 1.2955e-08 1.0000e-03 1.3005e-08 1.0000e-03
+ 1.3010e-08 0.0000e+00 1.3150e-08 0.0000e+00 1.3155e-08 1.0000e-03
+ 1.3205e-08 1.0000e-03 1.3210e-08 0.0000e+00 1.3750e-08 0.0000e+00
+ 1.3755e-08 1.0000e-03 1.3805e-08 1.0000e-03 1.3810e-08 0.0000e+00
+ 1.3950e-08 0.0000e+00 1.3955e-08 1.0000e-03 1.4005e-08 1.0000e-03
+ 1.4010e-08 0.0000e+00 1.4550e-08 0.0000e+00 1.4555e-08 1.0000e-03
+ 1.4605e-08 1.0000e-03 1.4610e-08 0.0000e+00 1.4750e-08 0.0000e+00
+ 1.4755e-08 1.0000e-03 1.4805e-08 1.0000e-03 1.4810e-08 0.0000e+00
+ 1.5350e-08 0.0000e+00 1.5355e-08 1.0000e-03 1.5405e-08 1.0000e-03
+ 1.5410e-08 0.0000e+00 1.5550e-08 0.0000e+00 1.5555e-08 1.0000e-03
+ 1.5605e-08 1.0000e-03 1.5610e-08 0.0000e+00 1.6150e-08 0.0000e+00
+ 1.6155e-08 1.0000e-03 1.6205e-08 1.0000e-03 1.6210e-08 0.0000e+00
+ 1.6350e-08 0.0000e+00 1.6355e-08 1.0000e-03 1.6405e-08 1.0000e-03
+ 1.6410e-08 0.0000e+00 1.6950e-08 0.0000e+00 1.6955e-08 1.0000e-03
+ 1.7005e-08 1.0000e-03 1.7010e-08 0.0000e+00 1.7150e-08 0.0000e+00
+ 1.7155e-08 1.0000e-03 1.7205e-08 1.0000e-03 1.7210e-08 0.0000e+00
+ 1.7750e-08 0.0000e+00 1.7755e-08 1.0000e-03 1.7805e-08 1.0000e-03
+ 1.7810e-08 0.0000e+00 1.7950e-08 0.0000e+00 1.7955e-08 1.0000e-03
+ 1.8005e-08 1.0000e-03 1.8010e-08 0.0000e+00 1.8550e-08 0.0000e+00
+ 1.8555e-08 1.0000e-03 1.8605e-08 1.0000e-03 1.8610e-08 0.0000e+00
+ 1.8750e-08 0.0000e+00 1.8755e-08 1.0000e-03 1.8805e-08 1.0000e-03
+ 1.8810e-08 0.0000e+00 1.9350e-08 0.0000e+00 1.9355e-08 1.0000e-03
+ 1.9405e-08 1.0000e-03 1.9410e-08 0.0000e+00 1.9550e-08 0.0000e+00
+ 1.9555e-08 1.0000e-03 1.9605e-08 1.0000e-03 1.9610e-08 0.0000e+00
+ 2.0150e-08 0.0000e+00 2.0155e-08 1.0000e-03 2.0205e-08 1.0000e-03
+ 2.0210e-08 0.0000e+00 2.0350e-08 0.0000e+00 2.0355e-08 1.0000e-03
+ 2.0405e-08 1.0000e-03 2.0410e-08 0.0000e+00 2.0950e-08 0.0000e+00
+ 2.0955e-08 1.0000e-03 2.1005e-08 1.0000e-03 2.1010e-08 0.0000e+00
+ 2.1150e-08 0.0000e+00 2.1155e-08 1.0000e-03 2.1205e-08 1.0000e-03
+ 2.1210e-08 0.0000e+00 2.1750e-08 0.0000e+00 2.1755e-08 1.0000e-03
+ 2.1805e-08 1.0000e-03 2.1810e-08 0.0000e+00 2.1950e-08 0.0000e+00
+ 2.1955e-08 1.0000e-03 2.2005e-08 1.0000e-03 2.2010e-08 0.0000e+00
+ 2.2550e-08 0.0000e+00 2.2555e-08 1.0000e-03 2.2605e-08 1.0000e-03
+ 2.2610e-08 0.0000e+00 2.2750e-08 0.0000e+00 2.2755e-08 1.0000e-03
+ 2.2805e-08 1.0000e-03 2.2810e-08 0.0000e+00 2.3350e-08 0.0000e+00
+ 2.3355e-08 1.0000e-03 2.3405e-08 1.0000e-03 2.3410e-08 0.0000e+00
+ 2.3550e-08 0.0000e+00 2.3555e-08 1.0000e-03 2.3605e-08 1.0000e-03
+ 2.3610e-08 0.0000e+00 2.4150e-08 0.0000e+00 2.4155e-08 1.0000e-03
+ 2.4205e-08 1.0000e-03 2.4210e-08 0.0000e+00 2.4350e-08 0.0000e+00
+ 2.4355e-08 1.0000e-03 2.4405e-08 1.0000e-03 2.4410e-08 0.0000e+00
+ 2.4950e-08 0.0000e+00 2.4955e-08 1.0000e-03 2.5005e-08 1.0000e-03
+ 2.5010e-08 0.0000e+00 2.5150e-08 0.0000e+00 2.5155e-08 1.0000e-03
+ 2.5205e-08 1.0000e-03 2.5210e-08 0.0000e+00 2.5750e-08 0.0000e+00
+ 2.5755e-08 1.0000e-03 2.5805e-08 1.0000e-03 2.5810e-08 0.0000e+00
+ 2.5950e-08 0.0000e+00 2.5955e-08 1.0000e-03 2.6005e-08 1.0000e-03
+ 2.6010e-08 0.0000e+00 2.6550e-08 0.0000e+00 2.6555e-08 1.0000e-03
+ 2.6605e-08 1.0000e-03 2.6610e-08 0.0000e+00 2.6750e-08 0.0000e+00
+ 2.6755e-08 1.0000e-03 2.6805e-08 1.0000e-03 2.6810e-08 0.0000e+00
+ 2.7350e-08 0.0000e+00 2.7355e-08 1.0000e-03 2.7405e-08 1.0000e-03
+ 2.7410e-08 0.0000e+00 2.7550e-08 0.0000e+00 2.7555e-08 1.0000e-03
+ 2.7605e-08 1.0000e-03 2.7610e-08 0.0000e+00 2.8150e-08 0.0000e+00
+ 2.8155e-08 1.0000e-03 2.8205e-08 1.0000e-03 2.8210e-08 0.0000e+00
+ 2.8350e-08 0.0000e+00 2.8355e-08 1.0000e-03 2.8405e-08 1.0000e-03
+ 2.8410e-08 0.0000e+00 2.8950e-08 0.0000e+00 2.8955e-08 1.0000e-03
+ 2.9005e-08 1.0000e-03 2.9010e-08 0.0000e+00 2.9150e-08 0.0000e+00
+ 2.9155e-08 1.0000e-03 2.9205e-08 1.0000e-03 2.9210e-08 0.0000e+00
+ 2.9750e-08 0.0000e+00 2.9755e-08 1.0000e-03 2.9805e-08 1.0000e-03
+ 2.9810e-08 0.0000e+00 2.9950e-08 0.0000e+00 2.9955e-08 1.0000e-03
+ 3.0005e-08 1.0000e-03 3.0010e-08 0.0000e+00 3.0550e-08 0.0000e+00
+ 3.0555e-08 1.0000e-03 3.0605e-08 1.0000e-03 3.0610e-08 0.0000e+00
+ 3.0750e-08 0.0000e+00 3.0755e-08 1.0000e-03 3.0805e-08 1.0000e-03
+ 3.0810e-08 0.0000e+00 3.1350e-08 0.0000e+00 3.1355e-08 1.0000e-03
+ 3.1405e-08 1.0000e-03 3.1410e-08 0.0000e+00 3.1550e-08 0.0000e+00
+ 3.1555e-08 1.0000e-03 3.1605e-08 1.0000e-03 3.1610e-08 0.0000e+00
+ 3.2150e-08 0.0000e+00 3.2155e-08 1.0000e-03 3.2205e-08 1.0000e-03
+ 3.2210e-08 0.0000e+00 3.2350e-08 0.0000e+00 3.2355e-08 1.0000e-03
+ 3.2405e-08 1.0000e-03 3.2410e-08 0.0000e+00)
IINBIAS1 0 INB11 pulse(0 0.001 550p 5p 5p 50p 200p)
ITARGET 0 TARGET0  PWL(0 0 20P 0 7.5000e-10 0.0000e+00 7.5500e-10 1.0000e-03 8.0500e-10 1.0000e-03
+ 8.1000e-10 0.0000e+00 9.5000e-10 0.0000e+00 9.5500e-10 1.0000e-03
+ 1.0050e-09 1.0000e-03 1.0100e-09 0.0000e+00 1.5500e-09 0.0000e+00
+ 1.5550e-09 1.0000e-03 1.6050e-09 1.0000e-03 1.6100e-09 0.0000e+00
+ 1.7500e-09 0.0000e+00 1.7550e-09 1.0000e-03 1.8050e-09 1.0000e-03
+ 1.8100e-09 0.0000e+00 2.3500e-09 0.0000e+00 2.3550e-09 1.0000e-03
+ 2.4050e-09 1.0000e-03 2.4100e-09 0.0000e+00 2.5500e-09 0.0000e+00
+ 2.5550e-09 1.0000e-03 2.6050e-09 1.0000e-03 2.6100e-09 0.0000e+00
+ 3.1500e-09 0.0000e+00 3.1550e-09 1.0000e-03 3.2050e-09 1.0000e-03
+ 3.2100e-09 0.0000e+00 3.3500e-09 0.0000e+00 3.3550e-09 1.0000e-03
+ 3.4050e-09 1.0000e-03 3.4100e-09 0.0000e+00 3.9500e-09 0.0000e+00
+ 3.9550e-09 1.0000e-03 4.0050e-09 1.0000e-03 4.0100e-09 0.0000e+00
+ 4.1500e-09 0.0000e+00 4.1550e-09 1.0000e-03 4.2050e-09 1.0000e-03
+ 4.2100e-09 0.0000e+00 4.7500e-09 0.0000e+00 4.7550e-09 1.0000e-03
+ 4.8050e-09 1.0000e-03 4.8100e-09 0.0000e+00 4.9500e-09 0.0000e+00
+ 4.9550e-09 1.0000e-03 5.0050e-09 1.0000e-03 5.0100e-09 0.0000e+00
+ 5.5500e-09 0.0000e+00 5.5550e-09 1.0000e-03 5.6050e-09 1.0000e-03
+ 5.6100e-09 0.0000e+00 5.7500e-09 0.0000e+00 5.7550e-09 1.0000e-03
+ 5.8050e-09 1.0000e-03 5.8100e-09 0.0000e+00 6.3500e-09 0.0000e+00
+ 6.3550e-09 1.0000e-03 6.4050e-09 1.0000e-03 6.4100e-09 0.0000e+00
+ 6.5500e-09 0.0000e+00 6.5550e-09 1.0000e-03 6.6050e-09 1.0000e-03
+ 6.6100e-09 0.0000e+00 7.1500e-09 0.0000e+00 7.1550e-09 1.0000e-03
+ 7.2050e-09 1.0000e-03 7.2100e-09 0.0000e+00 7.3500e-09 0.0000e+00
+ 7.3550e-09 1.0000e-03 7.4050e-09 1.0000e-03 7.4100e-09 0.0000e+00
+ 7.9500e-09 0.0000e+00 7.9550e-09 1.0000e-03 8.0050e-09 1.0000e-03
+ 8.0100e-09 0.0000e+00 8.1500e-09 0.0000e+00 8.1550e-09 1.0000e-03
+ 8.2050e-09 1.0000e-03 8.2100e-09 0.0000e+00 8.7500e-09 0.0000e+00
+ 8.7550e-09 1.0000e-03 8.8050e-09 1.0000e-03 8.8100e-09 0.0000e+00
+ 8.9500e-09 0.0000e+00 8.9550e-09 1.0000e-03 9.0050e-09 1.0000e-03
+ 9.0100e-09 0.0000e+00 9.5500e-09 0.0000e+00 9.5550e-09 1.0000e-03
+ 9.6050e-09 1.0000e-03 9.6100e-09 0.0000e+00 9.7500e-09 0.0000e+00
+ 9.7550e-09 1.0000e-03 9.8050e-09 1.0000e-03 9.8100e-09 0.0000e+00
+ 1.0350e-08 0.0000e+00 1.0355e-08 1.0000e-03 1.0405e-08 1.0000e-03
+ 1.0410e-08 0.0000e+00 1.0550e-08 0.0000e+00 1.0555e-08 1.0000e-03
+ 1.0605e-08 1.0000e-03 1.0610e-08 0.0000e+00 1.1150e-08 0.0000e+00
+ 1.1155e-08 1.0000e-03 1.1205e-08 1.0000e-03 1.1210e-08 0.0000e+00
+ 1.1350e-08 0.0000e+00 1.1355e-08 1.0000e-03 1.1405e-08 1.0000e-03
+ 1.1410e-08 0.0000e+00 1.1950e-08 0.0000e+00 1.1955e-08 1.0000e-03
+ 1.2005e-08 1.0000e-03 1.2010e-08 0.0000e+00 1.2150e-08 0.0000e+00
+ 1.2155e-08 1.0000e-03 1.2205e-08 1.0000e-03 1.2210e-08 0.0000e+00
+ 1.2750e-08 0.0000e+00 1.2755e-08 1.0000e-03 1.2805e-08 1.0000e-03
+ 1.2810e-08 0.0000e+00 1.2950e-08 0.0000e+00 1.2955e-08 1.0000e-03
+ 1.3005e-08 1.0000e-03 1.3010e-08 0.0000e+00 1.3550e-08 0.0000e+00
+ 1.3555e-08 1.0000e-03 1.3605e-08 1.0000e-03 1.3610e-08 0.0000e+00
+ 1.3750e-08 0.0000e+00 1.3755e-08 1.0000e-03 1.3805e-08 1.0000e-03
+ 1.3810e-08 0.0000e+00 1.4350e-08 0.0000e+00 1.4355e-08 1.0000e-03
+ 1.4405e-08 1.0000e-03 1.4410e-08 0.0000e+00 1.4550e-08 0.0000e+00
+ 1.4555e-08 1.0000e-03 1.4605e-08 1.0000e-03 1.4610e-08 0.0000e+00
+ 1.5150e-08 0.0000e+00 1.5155e-08 1.0000e-03 1.5205e-08 1.0000e-03
+ 1.5210e-08 0.0000e+00 1.5350e-08 0.0000e+00 1.5355e-08 1.0000e-03
+ 1.5405e-08 1.0000e-03 1.5410e-08 0.0000e+00 1.5950e-08 0.0000e+00
+ 1.5955e-08 1.0000e-03 1.6005e-08 1.0000e-03 1.6010e-08 0.0000e+00
+ 1.6150e-08 0.0000e+00 1.6155e-08 1.0000e-03 1.6205e-08 1.0000e-03
+ 1.6210e-08 0.0000e+00 1.6750e-08 0.0000e+00 1.6755e-08 1.0000e-03
+ 1.6805e-08 1.0000e-03 1.6810e-08 0.0000e+00 1.6950e-08 0.0000e+00
+ 1.6955e-08 1.0000e-03 1.7005e-08 1.0000e-03 1.7010e-08 0.0000e+00
+ 1.7550e-08 0.0000e+00 1.7555e-08 1.0000e-03 1.7605e-08 1.0000e-03
+ 1.7610e-08 0.0000e+00 1.7750e-08 0.0000e+00 1.7755e-08 1.0000e-03
+ 1.7805e-08 1.0000e-03 1.7810e-08 0.0000e+00 1.8350e-08 0.0000e+00
+ 1.8355e-08 1.0000e-03 1.8405e-08 1.0000e-03 1.8410e-08 0.0000e+00
+ 1.8550e-08 0.0000e+00 1.8555e-08 1.0000e-03 1.8605e-08 1.0000e-03
+ 1.8610e-08 0.0000e+00 1.9150e-08 0.0000e+00 1.9155e-08 1.0000e-03
+ 1.9205e-08 1.0000e-03 1.9210e-08 0.0000e+00 1.9350e-08 0.0000e+00
+ 1.9355e-08 1.0000e-03 1.9405e-08 1.0000e-03 1.9410e-08 0.0000e+00
+ 1.9950e-08 0.0000e+00 1.9955e-08 1.0000e-03 2.0005e-08 1.0000e-03
+ 2.0010e-08 0.0000e+00 2.0150e-08 0.0000e+00 2.0155e-08 1.0000e-03
+ 2.0205e-08 1.0000e-03 2.0210e-08 0.0000e+00 2.0750e-08 0.0000e+00
+ 2.0755e-08 1.0000e-03 2.0805e-08 1.0000e-03 2.0810e-08 0.0000e+00
+ 2.0950e-08 0.0000e+00 2.0955e-08 1.0000e-03 2.1005e-08 1.0000e-03
+ 2.1010e-08 0.0000e+00 2.1550e-08 0.0000e+00 2.1555e-08 1.0000e-03
+ 2.1605e-08 1.0000e-03 2.1610e-08 0.0000e+00 2.1750e-08 0.0000e+00
+ 2.1755e-08 1.0000e-03 2.1805e-08 1.0000e-03 2.1810e-08 0.0000e+00
+ 2.2350e-08 0.0000e+00 2.2355e-08 1.0000e-03 2.2405e-08 1.0000e-03
+ 2.2410e-08 0.0000e+00 2.2550e-08 0.0000e+00 2.2555e-08 1.0000e-03
+ 2.2605e-08 1.0000e-03 2.2610e-08 0.0000e+00 2.3150e-08 0.0000e+00
+ 2.3155e-08 1.0000e-03 2.3205e-08 1.0000e-03 2.3210e-08 0.0000e+00
+ 2.3350e-08 0.0000e+00 2.3355e-08 1.0000e-03 2.3405e-08 1.0000e-03
+ 2.3410e-08 0.0000e+00 2.3950e-08 0.0000e+00 2.3955e-08 1.0000e-03
+ 2.4005e-08 1.0000e-03 2.4010e-08 0.0000e+00 2.4150e-08 0.0000e+00
+ 2.4155e-08 1.0000e-03 2.4205e-08 1.0000e-03 2.4210e-08 0.0000e+00
+ 2.4750e-08 0.0000e+00 2.4755e-08 1.0000e-03 2.4805e-08 1.0000e-03
+ 2.4810e-08 0.0000e+00 2.4950e-08 0.0000e+00 2.4955e-08 1.0000e-03
+ 2.5005e-08 1.0000e-03 2.5010e-08 0.0000e+00 2.5550e-08 0.0000e+00
+ 2.5555e-08 1.0000e-03 2.5605e-08 1.0000e-03 2.5610e-08 0.0000e+00
+ 2.5750e-08 0.0000e+00 2.5755e-08 1.0000e-03 2.5805e-08 1.0000e-03
+ 2.5810e-08 0.0000e+00 2.6350e-08 0.0000e+00 2.6355e-08 1.0000e-03
+ 2.6405e-08 1.0000e-03 2.6410e-08 0.0000e+00 2.6550e-08 0.0000e+00
+ 2.6555e-08 1.0000e-03 2.6605e-08 1.0000e-03 2.6610e-08 0.0000e+00
+ 2.7150e-08 0.0000e+00 2.7155e-08 1.0000e-03 2.7205e-08 1.0000e-03
+ 2.7210e-08 0.0000e+00 2.7350e-08 0.0000e+00 2.7355e-08 1.0000e-03
+ 2.7405e-08 1.0000e-03 2.7410e-08 0.0000e+00 2.7950e-08 0.0000e+00
+ 2.7955e-08 1.0000e-03 2.8005e-08 1.0000e-03 2.8010e-08 0.0000e+00
+ 2.8150e-08 0.0000e+00 2.8155e-08 1.0000e-03 2.8205e-08 1.0000e-03
+ 2.8210e-08 0.0000e+00 2.8750e-08 0.0000e+00 2.8755e-08 1.0000e-03
+ 2.8805e-08 1.0000e-03 2.8810e-08 0.0000e+00 2.8950e-08 0.0000e+00
+ 2.8955e-08 1.0000e-03 2.9005e-08 1.0000e-03 2.9010e-08 0.0000e+00
+ 2.9550e-08 0.0000e+00 2.9555e-08 1.0000e-03 2.9605e-08 1.0000e-03
+ 2.9610e-08 0.0000e+00 2.9750e-08 0.0000e+00 2.9755e-08 1.0000e-03
+ 2.9805e-08 1.0000e-03 2.9810e-08 0.0000e+00 3.0350e-08 0.0000e+00
+ 3.0355e-08 1.0000e-03 3.0405e-08 1.0000e-03 3.0410e-08 0.0000e+00
+ 3.0550e-08 0.0000e+00 3.0555e-08 1.0000e-03 3.0605e-08 1.0000e-03
+ 3.0610e-08 0.0000e+00 3.1150e-08 0.0000e+00 3.1155e-08 1.0000e-03
+ 3.1205e-08 1.0000e-03 3.1210e-08 0.0000e+00 3.1350e-08 0.0000e+00
+ 3.1355e-08 1.0000e-03 3.1405e-08 1.0000e-03 3.1410e-08 0.0000e+00
+ 3.1950e-08 0.0000e+00 3.1955e-08 1.0000e-03 3.2005e-08 1.0000e-03
+ 3.2010e-08 0.0000e+00 3.2150e-08 0.0000e+00 3.2155e-08 1.0000e-03
+ 3.2205e-08 1.0000e-03 3.2210e-08 0.0000e+00)

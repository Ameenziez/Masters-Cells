#used to convert SFQ PULSE TO SHORT DC CURRENT PULSE
#EACH OF THESE ADDS 36 JJS...

.SUBCKT DCPULSER SFQIN CURRENTPULSEOUT

XSPLIT LSmitll_SPLITT SFQIN SFQ1 SFQ2
XJTL1 LSMITLL_JTLT SFQ1 SFQ1DELAYED
XJTL2 LSMITLL_JTLT SFQ1DELAYED SFQ1DELAYED2
XJTL3 LSMITLL_JTLT SFQ1DELAYED2 SFQ1DELAYED3
XMERGE LSMITLL_MERGET SFQ2 SFQ1DELAYED3 OUTPUT
XDC LSmitll_PTLRX_SFQDC OUTPUT CURRENTPULSEOUT

.ENDS DCPULSER
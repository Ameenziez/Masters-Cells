.subckt DELAY7 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R


XDELAY1 bfr B6 INPUT XIN1  DCIN DC6 0 DOUTRD1
XDELAY2 bfr A5 DOUTRD1 XIN2  DC6 DC7  0 DOUTRD2
XDELAY3 bfr B7 DOUTRD2 B6  DC8 DC7  0 DOUTRD3
XDELAY4 bfr A5 DOUTRD3 A6 DC8 DC9   0 DOUTRD4
XDELAY5 bfr B7 DOUTRD4 B8 DC10 DC9    0 DOUTRD5
XDELAY6 bfr XOUT2 DOUTRD5 A6 DC10 DC11  0 DOUTRD6
XDELAY7 bfrsplit2 XOUT1 DOUTRD6 B8 DCOUT DC11    OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R

.ENDS DELAY7
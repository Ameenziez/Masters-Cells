#file containing necessary components for neuron 

.subckt SYNAPSE DIN DOUTL DOUTR WEIGHTL WEIGHTR NODEM
#ISTORE 0 WEIGHTM PWL(0 0 20P -190U 3000p -190u 3001p -200u)
#ISTORE 0 WEIGHTM PWL(0 0 20P -10U)
LINPUT DIN 0 1p
LSTORE1 WEIGHTL NODEM 45.8p
LSTORE2 NODEM WEIGHTR 45.8p
KWEIGHT1 LWIN LSTORE1  -0.05
#KWEIGHT1 LWIN LSTORE1  -0.05
#UNCOMMENT SECOND COUPLING MAYBE...
#KWEIGHT2 LWIN LSTORE2 -0.05
#KWEIGHT3 LQ LSTORE1 -0.01
#KWEIGHT4 LQ LSTORE2 0.01
LWin 0 2  40p
L1 3 2 7p
L2 2 4 7p
RSHUNT1 3 0 0.07
RSHUNT2 4 0 0.07
B1 3 3par N1 jjmit area=0.5
B2 4 4par N2 jjmit area=0.5
LP1 3par 0 0.2p
LP2 4par 0 0.2p
LQ 2 0 40p
#rQ 2N 0 0.05
K1 L2 LINPUT -0.5
K2 LINPUT L1 -0.5
KOUT LQ LOUT 0.1
#koutoffset LOUT LSTORE1  0.01
LOUT DOUTL DOUTR 10p
.ends SYNAPSE

#FASTER
.subckt SYNAPSEfast DIN DOUTL DOUTR WEIGHTL WEIGHTR NODEM
#ISTORE 0 WEIGHTM PWL(0 0 20P -190U 3000p -190u 3001p -200u)
#ISTORE 0 WEIGHTM PWL(0 0 20P -10U)
LINPUT DIN 0 1p
LSTORE1 WEIGHTL NODEM 45.8p
LSTORE2 NODEM WEIGHTR 45.8p
KWEIGHT1 LWIN LSTORE1  -0.05
#KWEIGHT1 LWIN LSTORE1  -0.05
#UNCOMMENT SECOND COUPLING MAYBE...
#KWEIGHT2 LWIN LSTORE2 -0.05
#KWEIGHT3 LQ LSTORE1 -0.01
#KWEIGHT4 LQ LSTORE2 0.01
LWin 0 2  40p
L1 3 2 2p
L2 2 4 2p
RSHUNT1 3 0 0.5
RSHUNT2 4 0 0.5

B1 3 3par N1 jjmit area=0.5
B2 4 4par N2 jjmit area=0.5
LP1 3par 0 0.2p
LP2 4par 0 0.2p
LQ 2 0 20p
#rQ 2N 0 0.05
K1 L2  LINPUT -0.5
K2 LINPUT L1 -0.5
KOUT LQ LOUT 0.1
#koutoffset LOUT LSTORE1  0.01
LOUT DOUTL DOUTR 25p
.ends SYNAPSEfast


#fastest
.subckt SYNAPSEfastest DIN DOUTL DOUTR WEIGHTL WEIGHTR NODEM
LINPUT DIN 0 6.24p
LSTORE1 WEIGHTL NODEM 45.8p
LSTORE2 NODEM WEIGHTR 45.8p
KWEIGHT1 LWIN LSTORE1  -0.05
LWin 0 2  40p
L1 3 2 2p
L2 2 4 2p
RSHUNT1 3 0 1.4
RSHUNT2 4 0 1.4
B1 3 3par N1 jjmit area=0.5
B2 4 4par N2 jjmit area=0.5
LP1 3par 0 0.2p
LP2 4par 0 0.2p
LQ 2 0 20p
K1 L2  LINPUT -0.2
K2 LINPUT L1 -0.2
KOUT LQ LOUT -0.2
#WAS 35
LOUT DOUTL DOUTR 10P
#consider taking out lout but how do I couple then...
.ends SYNAPSEfastest







.subckt COMPARATOR DIN CLKIN CLKOUT DOUT 
#increase jj area to push saturation limit 1.1-1.2 works
#magnitude must be greater than 0.12
LCOMPX CLKIN CLKOUT 6p
KCOMP1 LCOMPX LCOMPL -0.233
KCOMP2 LCOMPR LCOMPX -0.233
LCOMPT DIN AMP3 1p
LCOMPL AMP4 AMP3 3p
LCOMPR AMP3 AMP5 3p
BCOMPL AMP4 0 AMP11 jjmit area=1.5
BCOMPR AMP5 0 AMP12 jjmit area=1.5
#was 3p
LCOMPQ AMP3 0 3p
LCOMPOUT DOUT 0 3.25p
KCOMPOUT LCOMPQ LCOMPOUT 0.2
#was 3p
#changed lq from 3P
.ends COMPARATOR






.subckt AQFP2RSFQ XIN XOUT AQFPIN RSFQOUT DCIN DCOUT
#EXCITATION CURRENT AND DC OFFSET INDUCTORS
LX XIN XOUT 15p
#WAS 6P CHANGED
#was 1.51p
LD DCIN DCOUT 6.51p
#MUTUAL INDUCATANCES
K1 LX LD 0.2322
K2 LX L1 -0.2284
K3 LD L1 -0.1559
K5 L2 LD 0.1559
K6 L2 LX 0.228
#FEED IN DATA 
#was 32.3p
LQ N0 AQFPIN 2.3p
L1 N1 N0  1.47p
L2 N2 N0  1.47p
B1 N1 P1 13 jjmit area=2
LP1 P1 0 0.2p
#was 1.6314
RSHUNT1 N1 0 0.6134
B2 N2 P2 14 jjmit area=2
LP2 P2 0 0.2p
RSHUNT2 N2 0 1.2
#using shunt of 1.2 works well
#RSHUNT2 N2 0 16.42
#commented shunt out bc it recommended it in paper
#WAS 0.6
Rif N2 JTL1 0.7
IB 0 JTL2 PWL(0 0 20ps 160u)
#WAS 123u had to increase to 150u
L3A JTL1 JTL2 2.7p
#WAS 2.4
L4A JTL2 JTL3 0.185p
#was 0.185
L5A JTL3 RSFQOUT 4.6p
#was 4.6
#was 5.33p
B3 JTL2 P3 15 jjmit area=1.39
LP3 P3 0 0.2p
RSHUNT3 JTL2 0 26.4
#was 26.4
B4 RSFQOUT P4 16 jjmit area=2.13
LP4 P4 0 0.2p
RSHUNT4 RSFQOUT 0 5.1
#was 5.1
#was 1.12 according to calcs but higher resistance gets higher Vout...
.ends AQFP2RSFQ




.subckt bfr XIN DIN XOUT DCIN DCOUT DOUTL DOUTR
B1 8 0 11 jjmit area=0.5
B2 9 0 12 jjmit area=0.5
#RSHUNT 8 0 10
#RSHUNT1 8 0 6
#RSHUNT2 9 0 6.7
K1 LX LD 0.2322
K2 LD LOUT 3.27E-5
K3 LX LOUT 3.68E-5
K4 LD LQ 4.9E-4
K5 LX LQ 5.11E-4
K6 LOUT LQ -0.3878
#was minus
K7 L2 LD -0.1556
K8 L2 LX -0.228
K9 LX L1 -0.2284
K10 LD L1 -0.1559
L1 8 7 1.51p
L2 7 9 1.51p
LD DCIN DCOUT 7.94p
LIN DIN 7 1.526p
#LOUT DOUTL DOUTR  10.3p
LOUT DOUTL DOUTR 5.3p
LQ 7 0 5.84p
#WAS 5.84P
LX XIN XOUT 6.51p
.ends bfr


.subckt bfrsplit2 XIN DIN XOUT DCIN DCOUT DOUTL1 DOUTR1 DOUTL2 DOUTR2 
B1 8 0 11 jjmit area=0.5
B2 9 0 12 jjmit area=0.5
K1 LX LD 0.2322
K2 LD LOUT1 3.27E-5
K3 LX LOUT1 3.68E-5
K4 LD LQ 4.9E-4
K5 LX LQ 5.11E-4
#K6 LOUT1 LQ -0.3878
K6 LOUT1 LQ -0.2878
#was minus
K7 L2 LD -0.1556
K8 L2 LX -0.228
K9 LX L1 -0.2284
K10 LD L1 -0.1559
K11 LD LOUT2 3.27E-5
K12 LX LOUT2 3.68E-5
#K13 LOUT2 LQ -0.3878
K13 LOUT2 LQ -0.2878
L1 8 7 1.51p
L2 7 9 1.51p
LD DCIN DCOUT 7.94p
LIN DIN 7 1.526p
#LOUT DOUTL DOUTR  10.3p
LOUT1 DOUTL1 DOUTR1 10.3p
LOUT2 DOUTL2 DOUTR2 10.3p
#can delete this one
LQ 7 0 28.84p
#WAS 5.84
LX XIN XOUT 6.51p

#RSHUNT2 9 0 4.9
.ends bfrsplit2

.subckt bfrsplit3 XIN DIN XOUT DCIN DCOUT DOUTL1 DOUTR1 DOUTL2 DOUTR2 DOUTL3 DOUTR3
B1 8 0 11 jjmit area=0.5
B2 9 0 12 jjmit area=0.5
K1 LX LD 0.2322
K2 LD LOUT1 3.27E-5
K3 LX LOUT1 3.68E-5
K4 LD LQ 4.9E-4
K5 LX LQ 5.11E-4
K6 LOUT1 LQ -0.3878
K7 L2 LD -0.1556
K8 L2 LX -0.228
K9 LX L1 -0.2284
K10 LD L1 -0.1559
K11 LD LOUT2 3.27E-5
K12 LX LOUT2 3.68E-5
K13 LOUT2 LQ -0.3878
K14 LD LOUT3 3.27E-5
K15 LX LOUT3 3.68E-5
K16 LOUT3 LQ -0.3878
L1 8 7 1.51p
L2 7 9 1.51p
LD DCIN DCOUT 7.94p
LIN DIN 7 1.526p
#RSHUNT2 9 0 7
#WAS 4.9
LOUT1 DOUTL1 DOUTR1 5.3p
LOUT2 DOUTL2 DOUTR2 5.3p
#can delete this one
LOUT3 DOUTL3 DOUTR3 5.3p
LQ 7 0 10.84p
#WAS 5.84
LX XIN XOUT 6.51p
.ends bfrsplit3


.subckt bfrsyn XIN DIN XOUT DCIN DCOUT DOUTL DOUTR
B1 8 0 11 jjmit area=0.5
B2 9 0 12 jjmit area=0.5
#RSHUNT 9 0 10
K1 LX LD 0.2322
K2 LD LOUT 3.27E-5
K3 LX LOUT 3.68E-5
K4 LD LQ 4.9E-4
K5 LX LQ 5.11E-4
K6 LOUT LQ -0.3878
#was minus
K7 L2 LD -0.1556
K8 L2 LX -0.228
K9 LX L1 -0.2284
K10 LD L1 -0.1559
L1 8 7 1.51p
L2 7 9 1.51p
LD DCIN DCOUT 7.94p
LIN DIN 7 1.526p
#LOUT DOUTL DOUTR  10.3p
LOUT DOUTL DOUTR 25.3p
LQ 7 0 30.84p
LX XIN XOUT 6.51p
.ends bfrsyn

.subckt bfrSHUNTED XIN DIN XOUT DCIN DCOUT DOUTL DOUTR
B1 8 0 11 jjmit area=0.5
B2 9 0 12 jjmit area=0.5
#RSHUNT 8 0 10
#RSHUNT1 8 0 6
RSHUNT2 9 0 4
K1 LX LD 0.2322
K2 LD LOUT 3.27E-5
K3 LX LOUT 3.68E-5
K4 LD LQ 4.9E-4
K5 LX LQ 5.11E-4
K6 LOUT LQ -0.3878
#was minus
K7 L2 LD -0.1556
K8 L2 LX -0.228
K9 LX L1 -0.2284
K10 LD L1 -0.1559
L1 8 7 1.51p
L2 7 9 1.51p
LD DCIN DCOUT 7.94p
LIN DIN 7 1.526p
#LOUT DOUTL DOUTR  10.3p
LOUT DOUTL DOUTR 20.3p
LQ 7 0 25.84p
#WAS 5.84P
LX XIN XOUT 6.51p
.ends bfr

.subckt bfrsplit4 XIN DIN XOUT DCIN DCOUT DOUTL1 DOUTR1 DOUTL2 DOUTR2 DOUTL3 DOUTR3 DOUTL4 DOUTR4
B1 8 0 11 jjmit area=0.5
B2 9 0 12 jjmit area=0.5
K1 LX LD 0.2322
K2 LD LOUT1 3.27E-5
K3 LX LOUT1 3.68E-5
K4 LD LQ 4.9E-4
K5 LX LQ 5.11E-4
K6 LOUT1 LQ -0.15878
K7 L2 LD -0.1556
K8 L2 LX -0.228
K9 LX L1 -0.2284
K10 LD L1 -0.1559
K11 LD LOUT2 3.27E-5
K12 LX LOUT2 3.68E-5
K13 LOUT2 LQ -0.15878
K14 LD LOUT3 3.27E-5
K15 LX LOUT3 3.68E-5
K16 LOUT3 LQ -0.15878
K17 LD LOUT4 3.27E-5
K18 LX LOUT4 3.68E-5
K19 LOUT4 LQ -0.15878
L1 8 7 1.51p
L2 7 9 1.51p
LD DCIN DCOUT 7.94p
LIN DIN 7 1.526p
#RSHUNT2 9 0 7
#WAS 6
LOUT1 DOUTL1 DOUTR1 10.3p
LOUT2 DOUTL2 DOUTR2 10.3p
#can delete this one
LOUT3 DOUTL3 DOUTR3 10.3p
LOUT4 DOUTL4 DOUTR4 10.3p
LQ 7 0 28.84p
#WAS 5.84
LX XIN XOUT 6.51p
.ends bfrsplit4


.subckt bfrconst XIN DIN XOUT DCIN DCOUT DOUTL DOUTR
B1 8 0 11 jjmit area=0.5
B2 9 0 12 jjmit area=0.5
#RSHUNT 8 0 10
#RSHUNT1 8 0 6
#RSHUNT2 9 0 6.7
K1 LX LD 0.2322
K2 LD LOUT 3.27E-5
K3 LX LOUT 3.68E-5
K4 LD LQ 4.9E-4
K5 LX LQ 5.11E-4
K6 LOUT LQ -0.3878
#was minus
K7 L2 LD -0.1556
K8 L2 LX -0.228
K9 LX L1 -0.2284
K10 LD L1 -0.1559
L1 8 7 1.51p
L2 7 9 1.51p
LD DCIN DCOUT 7.94p
LIN DIN 7 1.526p
#LOUT DOUTL DOUTR  10.3p
LOUT DOUTL DOUTR 25.3p
LQ 7 0 5.84p
#WAS 5.84P
LX XIN XOUT 6.51p
.ends bfrconst

.subckt bfrconst2 XIN DIN XOUT DCIN DCOUT DOUT1L DOUT1R DOUT2L DOUT2R
B1 8 0 11 jjmit area=0.5
B2 9 0 12 jjmit area=0.5
#RSHUNT 8 0 10
#RSHUNT1 8 0 6
#RSHUNT2 9 0 6.7
K1 LX LD 0.2322
K2 LD LOUT1 3.27E-5
K3 LX LOUT1 3.68E-5
K4 LD LQ 4.9E-4
K5 LX LQ 5.11E-4
K6 LOUT1 LQ -0.3878
K7 LOUT2 LQ -0.3878
K8 LD LOUT2 3.27E-5
K9 LX LOUT2 3.68E-5
#was minus
K7 L2 LD -0.1556
K8 L2 LX -0.228
K9 LX L1 -0.2284
K10 LD L1 -0.1559
L1 8 7 1.51p
L2 7 9 1.51p
LD DCIN DCOUT 7.94p
LIN DIN 7 1.526p
#LOUT DOUTL DOUTR  10.3p
LOUT1 DOUT1L DOUT1R 35.3p
LOUT2 DOUT2L DOUT2R 35.3p
LQ 7 0 25.84p
#WAS 5.84P
LX XIN XOUT 6.51p
.ends bfrconst2


.subckt bfrconv XIN DIN XOUT DCIN DCOUT DOUTL DOUTR
B1 8 0 11 jjmit area=0.5
B2 9 0 12 jjmit area=0.5
#RSHUNT 8 0 10
#RSHUNT1 8 0 6
#RSHUNT2 9 0 6.7
K1 LX LD 0.2322
K2 LD LOUT 3.27E-5
K3 LX LOUT 3.68E-5
K4 LD LQ 4.9E-4
K5 LX LQ 5.11E-4
K6 LOUT LQ -0.1178
#was 1.178
#0.1878
#WAS -0.3878
#was minus
K7 L2 LD -0.1556
K8 L2 LX -0.228
K9 LX L1 -0.2284
K10 LD L1 -0.1559
L1 8 7 1.51p
L2 7 9 1.51p
LD DCIN DCOUT 7.94p
LIN DIN 7 1.526p
#LOUT DOUTL DOUTR  10.3p
LOUT DOUTL DOUTR 20.3p
#WAS 25.3P
LQ 7 0 13.84p
#WAS 13.84
#WAS 5.84P
LX XIN XOUT 6.51p
.ends bfrconv



.subckt bfrsplit6 XIN DIN XOUT DCIN DCOUT DOUTL1 DOUTR1 DOUTL2 DOUTR2 DOUTL3 DOUTR3 DOUTL4 DOUTR4 DOUTL5 DOUTR5 DOUTL6 DOUTR6
B1 8 0 11 jjmit area=0.5
B2 9 0 12 jjmit area=0.5
K1 LX LD 0.2322
K2 LD LOUT1 3.27E-5
K3 LX LOUT1 3.68E-5
K4 LD LQ 4.9E-4
K5 LX LQ 5.11E-4
K6 LOUT1 LQ -0.10878
K7 L2 LD -0.1556
K8 L2 LX -0.228
K9 LX L1 -0.2284
K10 LD L1 -0.1559
K11 LD LOUT2 3.27E-5
K12 LX LOUT2 3.68E-5
K13 LOUT2 LQ -0.10878
K14 LD LOUT3 3.27E-5
K15 LX LOUT3 3.68E-5
K16 LOUT3 LQ -0.10878
K17 LD LOUT4 3.27E-5
K18 LX LOUT4 3.68E-5
K19 LOUT4 LQ -0.10878
K20 LD LOUT5 3.27E-5
K21 LX LOUT5 3.68E-5
K22 LOUT5 LQ -0.10878
K23 LD LOUT6 3.27E-5
K24 LX LOUT6 3.68E-5
K25 LOUT6 LQ -0.10878
L1 8 7 1.51p
L2 7 9 1.51p
LD DCIN DCOUT 7.94p
LIN DIN 7 1.526p
#WAS 6
LOUT1 DOUTL1 DOUTR1 10.3p
LOUT2 DOUTL2 DOUTR2 10.3p
#can delete this one
LOUT3 DOUTL3 DOUTR3 10.3p
LOUT4 DOUTL4 DOUTR4 10.3p
LOUT5 DOUTL5 DOUTR5 10.3p
LOUT6 DOUTL6 DOUTR6 10.3p
LQ 7 0 28.84p
#WAS 5.84
LX XIN XOUT 6.51p
.ends bfrsplit6


.model jjmit jj(rtype=1, vg=2.6m,
+ icrit=0.1m, r0=144, rn=16, cap=0.07p)
.ends componentsedit
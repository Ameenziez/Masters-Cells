
#works well!
#got the data to propagate
.include LSmitll_DCSFQ_PTLTX_v1p5.cir
.include LSmitll_bufft_v1p5.cir
.include LSmitll_PTLRX_SFQDC_v1p5.cir
.include LSmitll_SPLITT_v1p5.cir
.INCLUDE LSMITLL_JTLT_V1P5.CIR
.INCLUDE LSMITLL_MERGET_V1P5.CIR
.include storeedit.cir
.INCLUDE COMPONENTSEDIT.CIR
.INCLUDE COMP3.CIR
.INCLUDE COMP4.CIR
.INCLUDE COMP5.CIR
.INCLUDE COMP6.CIR
.include conv.cir
.INCLUDE synapsenext2.CIR
.INCLUDE DCPULSER.CIR
.INCLUDE MULTISPLIT.CIR
.include transmit.cir
.INCLUDE DELAY7.CIR
.INCLUDE AND.CIR
.INCLUDE AND3.CIR
.INCLUDE OR3.CIR
.include PERCEPTRON.CIR
.include PERCEPTRON2.CIR
.include CONVINTERFACE.cir


# TRY SHIFTING CLK OF OUTPUT BACK A BIT...

.tran 1ps 10000PS 0ps 1p
#MLP:
#D=Oi.T + Oi.!Oj + T.!Oj 

#setup circuitry
VAC1   A1   0   SIN(0 723mV 10GHz 200Ps 0)
RAC1   A1   A2   1000
LAC1   A2   A3   0.1p
VAC2   B1   0   SIN(0 723mV 10GHz 175.0ps 0)
RAC2   B1   B2   1000
LAC2   B2   B3   0.1p
VDC    DC1   0   pwl(0 0 20p 1023mV)
RDC    DC1   DC2   1000
LDC    DC2   DC3  0.1p
#VDCconv    DCc1   0   PWL(0ps 0mV 20ps 1023mV 1.881e-08 1023mV 1.8811000000000002e-08 0)
VDCconv    DCc1   0   PWL(0ps 0mV 20ps 1023mV)

RDCconv    DCc1   DCc2  640
LDCconv    DCc2   DCc3   0.1p




#SECOND LAYER SYNAPSE 1
IINITAL21 0 INITIAL21 PWL( 0 0 20P flx21*2*22.6U)
XSTORE21 BISTORE SFQOUTPLUS21 SFQOUTMINUS21 WEIGHTL21 WEIGHTR21


#NEXT LAYER BIAS
#Iactualsynbias21 0 ACTUALSYNB21x PWL(0 0 640P 0 665P 670U 700P 0 840P 0 865P 670U 900P 0  1040P 0 1065P 670U 1100P 0 1240P 0 1265P 670U 1300P 0  )
LSYNB21 ACTUALSYNB21x ACTUALSYNB21 1p  
KSYNB21 LSYNB21 LSYNADJUSTB21 0.3
LSYNADJUSTB21 0 ADJUSTB21 5P 

#SPLIT TARGET BETWEEN 2 NEURONS
LTARGET1 TARGET0 TARGET1 1p
LTARGET2 TARGET0 TARGET2 1p

#SPLIT INPUTS BETWEEN 2 NEURONS
LINPUT1 IN1 INPUT11 1P
#LINPUT2 IN1 INPUT12 1P
LINPUT3 IN2 INPUT13 1P
#LINPUT4 IN2 INPUT14 1P
LINPUTBIAS11 INB11 INPUTB12 1P
#LINPUTBIAS12 INB11 INPUTB13 1P
#LINPUTBIASTERM INPUTB13 0 0.1p

#LTERM2 INPUT12 0 6.5p
#LTERM4 INPUT14 0 6.5p
#LTERM5 INPUTB13 0 6.5P



IINITALB21 0 INITIALB21 PWL( 0 0 20P flxb21*2*-22.6U)
XSTOREB21 BISTORE SFQOUTPLUSB21 SFQOUTMINUSB21 WEIGHTLB21 WEIGHTRB21

X21 SYNAPSEfastestnext2 OUTPUTAXON DOUT22 DOUT21  WEIGHTL21 WEIGHTR21 INITIAL21
XB21 SYNAPSEfastestnext2 ACTUALSYNB21  0 DOUT22   WEIGHTLB21 WEIGHTRB21 INITIALB21

.param flx11 = 0
.param flx12 = 2
.param flx13 = 2
.param flx14 = 0
.param flxb11 = 1
.param flxb12 = -1
.param flx21 = -1
.param flx22 = 3
.param flxb21 = 0


IINITAL11 0 INITIAL11 PWL( 0 0 20P -22U*2*flx11)
IINITALB11 0 INITIALB11 PWL( 0 0 20P -22u*2*flxb11)
IINITAL13 0 INITIAL13 PWL( 0 0 20P -22U*2*flx13)


##FINAL ACTIVATION - this works 
ITHRESH11 0 THRESH11 PWL(0 0 20p 15U)
ITHRESH21 0 THRESH21 PWL(0 0 20p -5U)
#was like 23u
XACTfinal COMP6 A5 DOUT21 A6  DC6 DC5   DOUTFINAL1 0   DOUTFINAL2 0   DOUTFINAL3 0   DOUTFINAL4  0 DOUTFINAL5 0 DOUTFINAL6 0   THRESH21

XNEURON1 3NEURON2 INPUT11 INPUT13 INPUTB12 TARGET1 DOUTFINAL1 DOUTFINAL2 THRESH11 A3 A5 B3 B4 DC3 DC5 DCC3 DCC4  OUTPUT1 0    OUTPUT2 0 OUTPUTAXON DELAYEDTARGETP 0 0 DELAYEDTARGETN   DELAYEDTARGETP2 0   INITIAL11 INITIAL13 INITIALB11
          #x3NEURON2 INPUT1 INPUT2 INPUTBIAS TARGET DOUTFINAL1 DOUTFINAL2 THRESH XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT DCCIN DCCOUT OUTPUT OUTPUTAXON

xbfrout1 bfrsplit4 B4 DOUTFINAL3 B6 dc6 DC8  0 actfinaloutp actfinaloutn 0 0 actfinaloutp2  actfinaloutn2 0 


xtargetdelay bfr B6 DELAYEDTARGETp b6x dc8 dc8x delayedtargetp21 0
xtargetdelay2 bfr A6 delayedtargetp21 A6x dc8X dc8xx delayedtargetp22 0

XDELAYin DELAY10 OUTPUT1 b6x b6xx A6x A6xx DC8xx DC8xxx  0 DELAYin1   DELAYin2 0
#xinputdelay bfr a6x OUTPUT1 a6xx dc8xxx dc8xx  delayedinput0 0
#xinputdelay2 bfr b6x delayedinput0 b6xx dc8xxx dc8xxxx delayedinput1 0

#add more so same clk
#XPERCEPTRON21 PERCEPTRON   B6  B7 A7 A6   OUTPUT1  actfinaloutp actfinaloutn DELAYEDTARGETP   DC8 DC9 INCR21 DECR21
#XPERCEPTRON21 PERCEPTRON2LAYER2   B6  B7 A7 A6   OUTPUT1  actfinaloutp actfinaloutn DELAYEDTARGETP   DC8 DC9 INCR21 DECR21

XPERCEPTRON21 PERCEPTRON2LAYER2   b6xx  B7 A7 A6Xx   delayin1  actfinaloutp actfinaloutn delayedtargetp22   DC8xxx DC9 INCR21 DECR21

XCONVO CONV A7 A8   DCC5 DCC4  INCR21 DECR21 SFQOUTPLUS21 SFQOUTMINUS21

#XPERCEPTRONb21 PERCEPTRON   B7  B8 A9 A8   ADJUSTB21  actfinaloutp2 actfinaloutn2 DELAYEDTARGETP2   DC9 DC10 INCRb21 DECRb21
XPERCEPTRONb21 PERCEPTRON2LAYER   B7  0 A9 A8   ADJUSTB21  actfinaloutp2 actfinaloutn2 DELAYEDTARGETP2   DC9 0 INCRb21 DECRb21

XCONVb21 CONV A9 0   0 DCC5  INCRb21 DECRb21 SFQOUTPLUSb21 SFQOUTMINUSb21









.PRINT DEVII IIN1
.PRINT DEVII IIN2
.PRINT DEVII ITARGET
.PRINT PHASE LQ.XACT11.XNEURON1
.PRINT PHASE LQ.XACTfinal

.print phase lstore1.x11.XNEURON1
.print phase lstore1.x12.XNEURON1
.print phase lstore1.xb11.XNEURON1
.print phase lstore1.X21
.print phase lstore1.Xb21

#.PRINT PHASE LQ.XACTfinal




.SUBCKT 3NEURON2 INPUT1 INPUT2 INPUTBIAS TARGET ACTNEXT1 ACTNEXT2 THRESH XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT DCCIN DCCOUT OUTPUT1 OUTPUT1GND OUTPUT2 OUTPUT2GND OUTPUTAXON DELAYOUTTARGET3 DELAYOUTTARGET3GND DELAYOUTTARGET4 DELAYOUTTARGET4GND DELAYOUTTARGET5 DELAYOUTTARGET5GND INITIAL11 INITIAL12 INITIALB11

#INPUTS
LSYN11 INPUT1 SYN11 1p  
LSYN12 INPUT2 SYN12 1p  
LSYNB11 INPUTBIAS SYNB11 1p  
LTARGET1 TARGET TARGET1 1p
LTARGET2 TARGET1 0 1p

#COUPLINGS
KSYN11 LSYN11 LSYNADJUST11 -0.1
KSYN12 LSYN12 LSYNADJUST12 -0.1
KSYNB11 LSYNB11 LSYNADJUSTB11 -0.1
KT1 LTARGET1 LADJUSTTARGET1 -0.05
KT2 LTARGET2 LADJUSTTARGET2 -0.05
LSYNADJUST11 0 ADJUST11 5P 
LSYNADJUST12 0 ADJUST12 5P 
LSYNADJUSTB11 0 ADJUSTB11 5P 
LADJUSTTARGET1 0 ADJUSTTARGET1 5P
LADJUSTTARGET2 0 ADJUSTTARGET2 5P


#SYNAPSE 1
#IINITAL11 0 INITIAL11 PWL( 0 0 20P -80U)
XSTORE11 BISTORE SFQOUTPLUS11 SFQOUTMINUS11 WEIGHTL11 WEIGHTR11
X11 SYNAPSEfastest SYN11 DOUT12 DOUT11 WEIGHTL11 WEIGHTR11 INITIAL11
#l111 SFQOUTPLUS11 0 1p
#l112 SFQOUTMINUS11 0 1p

#SYNAPSE 2
#IINITAL12 0 INITIAL12 PWL( 0 0 20P -80U)
XSTORE12 BISTORE SFQOUTPLUS12 SFQOUTMINUS12 WEIGHTL12 WEIGHTR12
X12 SYNAPSEfastest SYN12 DOUT13 DOUT12 WEIGHTL12 WEIGHTR12 INITIAL12
#l121 SFQOUTPLUS12 0 1p
#l122 SFQOUTMINUSB12 0 1p

#SYNAPSE BIAS
#IINITALB11 0 INITIALB11 PWL( 0 0 20P -80U)
XSTOREB11 BISTORE SFQOUTPLUSB11 SFQOUTMINUSB11 WEIGHTLB11 WEIGHTRB11
XB11 SYNAPSEfastest SYNB11 0 DOUT13 WEIGHTLB11 WEIGHTRB11 INITIALB11
#lB111 SFQOUTPLUSB11 0 1p
#lB112 SFQOUTMINUSB11 0 1p

#ACTIVATION
XACT11 COMP5 XIN1 DOUT11 A4 DCIN DC4 DOUTL11 0  0 DOUTR12  0 DOUTL13 OUTPUT1GND OUTPUT1 OUTPUT2GND OUTPUT2   THRESH

#AXON FOR OUTPUT
XTRANSMIT1 TRANSMIT DOUTL11 XIN2 B4 A4 A6 DC4 DC6 DCCIN DCC4 OUTPUTAXON

#DELAYS
XDELAYACT1 DELAY10 DOUTR12 B4 B5 A6 A7 DC6 DC7  DELAYOUT1 0  DELAYOUT2 0
XDELAYTARGET DELAY14 ADJUSTTARGET1 B5 B6 A7 A8 DC7 DC8  DELAYOUTTARGET1  0 DELAYOUTTARGET2 0
#XDELAYTARGET2 DELAY103 ADJUSTTARGET2 B7 B8 A9 A10 DC9 DC10  DELAYOUTTARGET3 DELAYOUTTARGET3GND   DELAYOUTTARGET4 DELAYOUTTARGET4GND DELAYOUTTARGET5  DELAYOUTTARGET5GND 
XDELAYTARGET2 DELAY143 ADJUSTTARGET2 B7 B8 A9 A10 DC9 DC10  DELAYOUTTARGET3 DELAYOUTTARGET3GND   DELAYOUTTARGET4 DELAYOUTTARGET4GND DELAYOUTTARGET5  DELAYOUTTARGET5GND 
#i think this was delay143


#LEARNING ALGORITHMS
#ASSUME DOUTFINAL1 0 DOUTFINAL2 0  DOUTFINAL3 0  0 DOUTFINAL4
#XMLP MLPNEW B6 B7 A8 A9 DELAYOUT1 DELAYOUT2 DELAYOUTTARGET1 DELAYOUTTARGET2 ACTNEXT1 ACTNEXT2 DC8 DC9 OUTPUTTARGET1L 0 OUTPUTTARGET2L 0 OUTPUTTARGET3L 0
#XDELAYTARGET2 DELAY18 ADJUSTTARGET2 B7 B8 A9 A10 DC9 dc10  DELAYOUTTARGET3GND DELAYOUTTARGET3  DELAYOUTTARGET4 DELAYOUTTARGET4GND  DELAYOUTTARGET5GND DELAYOUTTARGET5 
XMLP MLPNEW B6 B7 A8 A9 DELAYOUT1 DELAYOUT2 DELAYOUTTARGET1 DELAYOUTTARGET2 ACTNEXT1 ACTNEXT2 DC8 DC9   OUTPUTTARGET1L 0 OUTPUTTARGET2L 0 OUTPUTTARGET3L 0

XDELAYINPUT1 DELAY18 ADJUST11  B8  B9  A10 A11 DC10 DC11 DELAYOUTINPUT111 0 DELAYOUTINPUT112 0 DELAYOUTINPUT113 0 DELAYOUTINPUT114 0 DELAYOUTINPUT115 0 DELAYOUTINPUT116 0
XDELAYINPUT2 DELAY18 ADJUST12  B9  B10  A11 A12 DC11 DC12 DELAYOUTINPUT121 0 DELAYOUTINPUT122 0 DELAYOUTINPUT123 0 DELAYOUTINPUT124 0 DELAYOUTINPUT125 0 DELAYOUTINPUT126 0
XDELAYINPUTB1 DELAY18 ADJUSTB11  B10  B11  A12 A13 DC12 DC13 DELAYOUTINPUT1B1 0 DELAYOUTINPUT1B2 0 DELAYOUTINPUT1B3 0 DELAYOUTINPUT1B4 0 DELAYOUTINPUT1B5 0 DELAYOUTINPUT1B6 0

XDELAYact2 DELAY15 DOUTL13  B11 B12  A13 A14 DC13 DC14  DELAYOUTact111 0 0  DELAYOUTact112 DELAYOUTact113 0 0  DELAYOUTact114   DELAYOUTact115  0 0  DELAYOUTact116 
#XDELAYact2 DELAY15 DOUTL13  B11 B12  A13 A14 DC13 DC14  0 DELAYOUTact111 DELAYOUTact112 0 DELAYOUTact113 0 0  DELAYOUTact114   DELAYOUTact115  0 0  DELAYOUTact116 


XPERCEPTRON11 PERCEPTRON  B13 B12  A14 A15  DELAYOUTINPUT111 DELAYOUTact111 DELAYOUTact112 OUTPUTTARGET1L DC15 DC14 INCR11 DECR11
XPERCEPTRON12 PERCEPTRON  B14 B13  A15 A16  DELAYOUTINPUT121 DELAYOUTact113 DELAYOUTact114 OUTPUTTARGET2L DC16 DC15 INCR12 DECR12
XPERCEPTRONB11 PERCEPTRON  XOUT2 B14  A16 A17  DELAYOUTINPUT1B1 DELAYOUTact115 DELAYOUTact116 OUTPUTTARGET3L DCOUT DC16 INCRB11 DECRB11

XCONV11 CONV A17 A18 DCC5 DCC4 INCR11 DECR11 SFQOUTPLUS11 SFQOUTMINUS11
XCONV12 CONV A18 A19 DCC6 DCC5 INCR12 DECR12 SFQOUTPLUS12 SFQOUTMINUS12
XCONVB11 CONV A19 XOUT1 DCCOUT DCC6 INCRB11 DECRB11 SFQOUTPLUSB11 SFQOUTMINUSB11

.ENDS 3NEURON2


.SUBCKT MLPNEW XIN1 XOUT1 XIN2 XOUT2 OI1 OI2 T1 T2 OJ1 OJ2 DCIN DCOUT OUTPUTTARGET1L OUTPUTTARGET1R OUTPUTTARGET2L OUTPUTTARGET2R OUTPUTTARGET3L OUTPUTTARGET3R
#Oi.T
Xand1  AND  B7 XIN1  XIN2 A9  OI1 T1 DC9 DCIN  andout1
#Oi.!Oj
Xand2  AND B8 B7 A9 A10 OI2 OJ1 DC10 DC9 andout2
#T.!Oj
Xand3  AND B9 B8 A10 A11 T2 OJ2 DC11 DC10 andout3
#D=Oi.T + Oi.!Oj + T.!Oj 
X3OR OR3 B9 XOUT1 XOUT2 A11   ANDOUT1 ANDOUT2 ANDOUT3 DCOUT DC11  OUTPUTTARGET1L OUTPUTTARGET1R OUTPUTTARGET2L OUTPUTTARGET2R OUTPUTTARGET3L OUTPUTTARGET3R 
.ENDS MLPNEW













.SUBCKT DELAY10 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 XOUT1  DC15 DC14      DELAYOUT9 0
XDELAY10 bfrsplit2 XOUT2 DELAYOUT9 A10   DC15 DCOUT      OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R
.ends DELAY10


.SUBCKT DELAY103 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R  OUTPUT3L OUTPUT3R

XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR XOUT2 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 bfrsplit3 XOUT1 DELAYOUT6 B7  DCOUT DC12 OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R

.ends DELAY103


.SUBCKT DELAY11 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR XOUT2 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 bfrsplit2 XOUT1 DELAYOUT10 B9   DCOUT DC16   OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R

.ends DELAY11


.SUBCKT DELAY113 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR XOUT2 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 bfrsplit3 XOUT1 DELAYOUT10 B9   DCOUT DC16   OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R

.ends DELAY113




.SUBCKT DELAY14 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R

XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR A11 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 BFR B10 DELAYOUT10 B9   DC17 DC16   DELAYOUT11 0
XDELAY12 BFR A11 DELAYOUT11 A12   DC17 DC18  DELAYOUT12 0
XDELAY13 BFR B10 DELAYOUT12 XOUT1  DC19 DC18  DELAYOUT13 0
XDELAY14 bfrsplit2 XOUT2 DELAYOUT13 A12  DC19 DCOUT  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R
#XDELAY14 bfrsplit5 XOUT2 DELAYOUT13 A12  DC19 DCOUT  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R OUTPUT4L OUTPUT4R OUTPUT5L OUTPUT5R

.ends DELAY14


.SUBCKT DELAY143 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R

XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR A11 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 BFR B10 DELAYOUT10 B9   DC17 DC16   DELAYOUT11 0
XDELAY12 BFR A11 DELAYOUT11 A12   DC17 DC18  DELAYOUT12 0
XDELAY13 BFR B10 DELAYOUT12 XOUT1  DC19 DC18  DELAYOUT13 0
XDELAY14 bfrsplit3 XOUT2 DELAYOUT13 A12  DC19 DCOUT  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R
#XDELAY14 bfrsplit5 XOUT2 DELAYOUT13 A12  DC19 DCOUT  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R OUTPUT4L OUTPUT4R OUTPUT5L OUTPUT5R

.ends DELAY143

.SUBCKT DELAY15 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R OUTPUT4L OUTPUT4R OUTPUT5L OUTPUT5R OUTPUT6L OUTPUT6R
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR A11 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 BFR B10 DELAYOUT10 B9   DC17 DC16   DELAYOUT11 0
XDELAY12 BFR A11 DELAYOUT11 A12   DC17 DC18  DELAYOUT12 0
XDELAY13 BFR B10 DELAYOUT12 B11  DC19 DC18  DELAYOUT13 0
XDELAY14 BFR XOUT2 DELAYOUT13 A12  DC19 DC20  DELAYOUT14 0

XDELAY15 bfrsplit6 XOUT1 DELAYOUT14 B11 DCOUT DC20  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R OUTPUT4L OUTPUT4R OUTPUT5L OUTPUT5R OUTPUT6L OUTPUT6R

.ends DELAY15

.SUBCKT DELAY153 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R 
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR A11 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 BFR B10 DELAYOUT10 B9   DC17 DC16   DELAYOUT11 0
XDELAY12 BFR A11 DELAYOUT11 A12   DC17 DC18  DELAYOUT12 0
XDELAY13 BFR B10 DELAYOUT12 B11  DC19 DC18  DELAYOUT13 0
XDELAY14 BFR XOUT2 DELAYOUT13 A12  DC19 DC20  DELAYOUT14 0

XDELAY15 bfrsplit3 XOUT1 DELAYOUT14 B11 DCOUT DC20  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R 

.ends DELAY153



.SUBCKT DELAY16 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR A11 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 BFR B10 DELAYOUT10 B9   DC17 DC16   DELAYOUT11 0
XDELAY12 BFR A11 DELAYOUT11 A12   DC17 DC18  DELAYOUT12 0
XDELAY13 BFR B10 DELAYOUT12 B11  DC19 DC18  DELAYOUT13 0
XDELAY14 BFR A13 DELAYOUT13 A12  DC19 DC20  DELAYOUT14 0
XDELAY15 BFR XOUT1 DELAYOUT14 B11  DC21 DC20  DELAYOUT15 0
XDELAY16 bfrsplit2 A13 DELAYOUT15 XOUT2  DC21 DCOUT  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R
.ends DELAY16

.SUBCKT DELAY163 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR A11 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 BFR B10 DELAYOUT10 B9   DC17 DC16   DELAYOUT11 0
XDELAY12 BFR A11 DELAYOUT11 A12   DC17 DC18  DELAYOUT12 0
XDELAY13 BFR B10 DELAYOUT12 B11  DC19 DC18  DELAYOUT13 0
XDELAY14 BFR A13 DELAYOUT13 A12  DC19 DC20  DELAYOUT14 0
XDELAY15 BFR XOUT1 DELAYOUT14 B11  DC21 DC20  DELAYOUT15 0
XDELAY16 bfrsplit3 A13 DELAYOUT15 XOUT2  DC21 DCOUT  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R
.ends DELAY163


.SUBCKT DELAY18 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR A11 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 BFR B10 DELAYOUT10 B9   DC17 DC16   DELAYOUT11 0
XDELAY12 BFR A11 DELAYOUT11 A12   DC17 DC18  DELAYOUT12 0
XDELAY13 BFR B10 DELAYOUT12 B11  DC19 DC18  DELAYOUT13 0
XDELAY14 BFR A13 DELAYOUT13 A12  DC19 DC20  DELAYOUT14 0
XDELAY15 BFR B12 DELAYOUT14 B11  DC21 DC20  DELAYOUT15 0
XDELAY16 BFR A13 DELAYOUT15 A14  DC21 DC22  DELAYOUT16 0
XDELAY17 BFR B12 DELAYOUT16 XOUT1  DC23 DC22  DELAYOUT17 0
XDELAY18 bfrsplit3 XOUT2 DELAYOUT17 A14 DC23 DCOUT  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R  OUTPUT3L OUTPUT3R


.ends DELAY18

***    INPUTS  ***
IIN1 0 IN1 PWL(0 0 20P 0 1.55000e-09 0.00000e+00 1.55500e-09 1.00000e-03 1.60500e-09 1.00000e-03
+ 1.61000e-09 0.00000e+00 3.55000e-09 0.00000e+00 3.55500e-09 1.00000e-03
+ 3.60500e-09 1.00000e-03 3.61000e-09 0.00000e+00 5.55000e-09 0.00000e+00
+ 5.55500e-09 1.00000e-03 5.60500e-09 1.00000e-03 5.61000e-09 0.00000e+00
+ 7.55000e-09 0.00000e+00 7.55500e-09 1.00000e-03 7.60500e-09 1.00000e-03
+ 7.61000e-09 0.00000e+00 9.55000e-09 0.00000e+00 9.55500e-09 1.00000e-03
+ 9.60500e-09 1.00000e-03 9.61000e-09 0.00000e+00 1.15500e-08 0.00000e+00
+ 1.15550e-08 1.00000e-03 1.16050e-08 1.00000e-03 1.16100e-08 0.00000e+00
+ 1.35500e-08 0.00000e+00 1.35550e-08 1.00000e-03 1.36050e-08 1.00000e-03
+ 1.36100e-08 0.00000e+00 1.55500e-08 0.00000e+00 1.55550e-08 1.00000e-03
+ 1.56050e-08 1.00000e-03 1.56100e-08 0.00000e+00 1.75500e-08 0.00000e+00
+ 1.75550e-08 1.00000e-03 1.76050e-08 1.00000e-03 1.76100e-08 0.00000e+00
+ 1.95500e-08 0.00000e+00 1.95550e-08 1.00000e-03 1.96050e-08 1.00000e-03
+ 1.96100e-08 0.00000e+00 2.15500e-08 0.00000e+00 2.15550e-08 1.00000e-03
+ 2.16050e-08 1.00000e-03 2.16100e-08 0.00000e+00 2.35500e-08 0.00000e+00
+ 2.35550e-08 1.00000e-03 2.36050e-08 1.00000e-03 2.36100e-08 0.00000e+00
+ 2.55500e-08 0.00000e+00 2.55550e-08 1.00000e-03 2.56050e-08 1.00000e-03
+ 2.56100e-08 0.00000e+00 2.75500e-08 0.00000e+00 2.75550e-08 1.00000e-03
+ 2.76050e-08 1.00000e-03 2.76100e-08 0.00000e+00 2.95500e-08 0.00000e+00
+ 2.95550e-08 1.00000e-03 2.96050e-08 1.00000e-03 2.96100e-08 0.00000e+00
+ 3.15500e-08 0.00000e+00 3.15550e-08 1.00000e-03 3.16050e-08 1.00000e-03
+ 3.16100e-08 0.00000e+00 3.35500e-08 0.00000e+00 3.35550e-08 1.00000e-03
+ 3.36050e-08 1.00000e-03 3.36100e-08 0.00000e+00 3.55500e-08 0.00000e+00
+ 3.55550e-08 1.00000e-03 3.56050e-08 1.00000e-03 3.56100e-08 0.00000e+00
+ 3.75500e-08 0.00000e+00 3.75550e-08 1.00000e-03 3.76050e-08 1.00000e-03
+ 3.76100e-08 0.00000e+00 3.95500e-08 0.00000e+00 3.95550e-08 1.00000e-03
+ 3.96050e-08 1.00000e-03 3.96100e-08 0.00000e+00 4.15500e-08 0.00000e+00
+ 4.15550e-08 1.00000e-03 4.16050e-08 1.00000e-03 4.16100e-08 0.00000e+00
+ 4.35500e-08 0.00000e+00 4.35550e-08 1.00000e-03 4.36050e-08 1.00000e-03
+ 4.36100e-08 0.00000e+00 4.55500e-08 0.00000e+00 4.55550e-08 1.00000e-03
+ 4.56050e-08 1.00000e-03 4.56100e-08 0.00000e+00 4.75500e-08 0.00000e+00
+ 4.75550e-08 1.00000e-03 4.76050e-08 1.00000e-03 4.76100e-08 0.00000e+00
+ 4.95500e-08 0.00000e+00 4.95550e-08 1.00000e-03 4.96050e-08 1.00000e-03
+ 4.96100e-08 0.00000e+00 5.15500e-08 0.00000e+00 5.15550e-08 1.00000e-03
+ 5.16050e-08 1.00000e-03 5.16100e-08 0.00000e+00 5.35500e-08 0.00000e+00
+ 5.35550e-08 1.00000e-03 5.36050e-08 1.00000e-03 5.36100e-08 0.00000e+00
+ 5.55500e-08 0.00000e+00 5.55550e-08 1.00000e-03 5.56050e-08 1.00000e-03
+ 5.56100e-08 0.00000e+00 5.75500e-08 0.00000e+00 5.75550e-08 1.00000e-03
+ 5.76050e-08 1.00000e-03 5.76100e-08 0.00000e+00 5.95500e-08 0.00000e+00
+ 5.95550e-08 1.00000e-03 5.96050e-08 1.00000e-03 5.96100e-08 0.00000e+00
+ 6.15500e-08 0.00000e+00 6.15550e-08 1.00000e-03 6.16050e-08 1.00000e-03
+ 6.16100e-08 0.00000e+00 6.35500e-08 0.00000e+00 6.35550e-08 1.00000e-03
+ 6.36050e-08 1.00000e-03 6.36100e-08 0.00000e+00 6.55500e-08 0.00000e+00
+ 6.55550e-08 1.00000e-03 6.56050e-08 1.00000e-03 6.56100e-08 0.00000e+00
+ 6.75500e-08 0.00000e+00 6.75550e-08 1.00000e-03 6.76050e-08 1.00000e-03
+ 6.76100e-08 0.00000e+00 6.95500e-08 0.00000e+00 6.95550e-08 1.00000e-03
+ 6.96050e-08 1.00000e-03 6.96100e-08 0.00000e+00 7.15500e-08 0.00000e+00
+ 7.15550e-08 1.00000e-03 7.16050e-08 1.00000e-03 7.16100e-08 0.00000e+00
+ 7.35500e-08 0.00000e+00 7.35550e-08 1.00000e-03 7.36050e-08 1.00000e-03
+ 7.36100e-08 0.00000e+00 7.55500e-08 0.00000e+00 7.55550e-08 1.00000e-03
+ 7.56050e-08 1.00000e-03 7.56100e-08 0.00000e+00 7.75500e-08 0.00000e+00
+ 7.75550e-08 1.00000e-03 7.76050e-08 1.00000e-03 7.76100e-08 0.00000e+00
+ 7.95500e-08 0.00000e+00 7.95550e-08 1.00000e-03 7.96050e-08 1.00000e-03
+ 7.96100e-08 0.00000e+00 8.15500e-08 0.00000e+00 8.15550e-08 1.00000e-03
+ 8.16050e-08 1.00000e-03 8.16100e-08 0.00000e+00 8.35500e-08 0.00000e+00
+ 8.35550e-08 1.00000e-03 8.36050e-08 1.00000e-03 8.36100e-08 0.00000e+00
+ 8.55500e-08 0.00000e+00 8.55550e-08 1.00000e-03 8.56050e-08 1.00000e-03
+ 8.56100e-08 0.00000e+00 8.75500e-08 0.00000e+00 8.75550e-08 1.00000e-03
+ 8.76050e-08 1.00000e-03 8.76100e-08 0.00000e+00 8.95500e-08 0.00000e+00
+ 8.95550e-08 1.00000e-03 8.96050e-08 1.00000e-03 8.96100e-08 0.00000e+00
+ 9.15500e-08 0.00000e+00 9.15550e-08 1.00000e-03 9.16050e-08 1.00000e-03
+ 9.16100e-08 0.00000e+00 9.35500e-08 0.00000e+00 9.35550e-08 1.00000e-03
+ 9.36050e-08 1.00000e-03 9.36100e-08 0.00000e+00 9.55500e-08 0.00000e+00
+ 9.55550e-08 1.00000e-03 9.56050e-08 1.00000e-03 9.56100e-08 0.00000e+00
+ 9.75500e-08 0.00000e+00 9.75550e-08 1.00000e-03 9.76050e-08 1.00000e-03
+ 9.76100e-08 0.00000e+00 9.95500e-08 0.00000e+00 9.95550e-08 1.00000e-03
+ 9.96050e-08 1.00000e-03 9.96100e-08 0.00000e+00 1.01550e-07 0.00000e+00
+ 1.01555e-07 1.00000e-03 1.01605e-07 1.00000e-03 1.01610e-07 0.00000e+00
+ 1.03550e-07 0.00000e+00 1.03555e-07 1.00000e-03 1.03605e-07 1.00000e-03
+ 1.03610e-07 0.00000e+00 1.05550e-07 0.00000e+00 1.05555e-07 1.00000e-03
+ 1.05605e-07 1.00000e-03 1.05610e-07 0.00000e+00 1.07550e-07 0.00000e+00
+ 1.07555e-07 1.00000e-03 1.07605e-07 1.00000e-03 1.07610e-07 0.00000e+00
+ 1.09550e-07 0.00000e+00 1.09555e-07 1.00000e-03 1.09605e-07 1.00000e-03
+ 1.09610e-07 0.00000e+00 1.11550e-07 0.00000e+00 1.11555e-07 1.00000e-03
+ 1.11605e-07 1.00000e-03 1.11610e-07 0.00000e+00 1.13550e-07 0.00000e+00
+ 1.13555e-07 1.00000e-03 1.13605e-07 1.00000e-03 1.13610e-07 0.00000e+00
+ 1.15550e-07 0.00000e+00 1.15555e-07 1.00000e-03 1.15605e-07 1.00000e-03
+ 1.15610e-07 0.00000e+00 1.17550e-07 0.00000e+00 1.17555e-07 1.00000e-03
+ 1.17605e-07 1.00000e-03 1.17610e-07 0.00000e+00 1.19550e-07 0.00000e+00
+ 1.19555e-07 1.00000e-03 1.19605e-07 1.00000e-03 1.19610e-07 0.00000e+00
+ 1.21550e-07 0.00000e+00 1.21555e-07 1.00000e-03 1.21605e-07 1.00000e-03
+ 1.21610e-07 0.00000e+00 1.23550e-07 0.00000e+00 1.23555e-07 1.00000e-03
+ 1.23605e-07 1.00000e-03 1.23610e-07 0.00000e+00 1.25550e-07 0.00000e+00
+ 1.25555e-07 1.00000e-03 1.25605e-07 1.00000e-03 1.25610e-07 0.00000e+00
+ 1.27550e-07 0.00000e+00 1.27555e-07 1.00000e-03 1.27605e-07 1.00000e-03
+ 1.27610e-07 0.00000e+00 1.29550e-07 0.00000e+00 1.29555e-07 1.00000e-03
+ 1.29605e-07 1.00000e-03 1.29610e-07 0.00000e+00 1.31550e-07 0.00000e+00
+ 1.31555e-07 1.00000e-03 1.31605e-07 1.00000e-03 1.31610e-07 0.00000e+00
+ 1.33550e-07 0.00000e+00 1.33555e-07 1.00000e-03 1.33605e-07 1.00000e-03
+ 1.33610e-07 0.00000e+00 1.35550e-07 0.00000e+00 1.35555e-07 1.00000e-03
+ 1.35605e-07 1.00000e-03 1.35610e-07 0.00000e+00 1.37550e-07 0.00000e+00
+ 1.37555e-07 1.00000e-03 1.37605e-07 1.00000e-03 1.37610e-07 0.00000e+00
+ 1.39550e-07 0.00000e+00 1.39555e-07 1.00000e-03 1.39605e-07 1.00000e-03
+ 1.39610e-07 0.00000e+00 1.41550e-07 0.00000e+00 1.41555e-07 1.00000e-03
+ 1.41605e-07 1.00000e-03 1.41610e-07 0.00000e+00 1.43550e-07 0.00000e+00
+ 1.43555e-07 1.00000e-03 1.43605e-07 1.00000e-03 1.43610e-07 0.00000e+00
+ 1.45550e-07 0.00000e+00 1.45555e-07 1.00000e-03 1.45605e-07 1.00000e-03
+ 1.45610e-07 0.00000e+00 1.47550e-07 0.00000e+00 1.47555e-07 1.00000e-03
+ 1.47605e-07 1.00000e-03 1.47610e-07 0.00000e+00 1.49550e-07 0.00000e+00
+ 1.49555e-07 1.00000e-03 1.49605e-07 1.00000e-03 1.49610e-07 0.00000e+00
+ 1.51550e-07 0.00000e+00 1.51555e-07 1.00000e-03 1.51605e-07 1.00000e-03
+ 1.51610e-07 0.00000e+00 1.53550e-07 0.00000e+00 1.53555e-07 1.00000e-03
+ 1.53605e-07 1.00000e-03 1.53610e-07 0.00000e+00 1.55550e-07 0.00000e+00
+ 1.55555e-07 1.00000e-03 1.55605e-07 1.00000e-03 1.55610e-07 0.00000e+00
+ 1.57550e-07 0.00000e+00 1.57555e-07 1.00000e-03 1.57605e-07 1.00000e-03
+ 1.57610e-07 0.00000e+00 1.59550e-07 0.00000e+00 1.59555e-07 1.00000e-03
+ 1.59605e-07 1.00000e-03 1.59610e-07 0.00000e+00 1.61550e-07 0.00000e+00
+ 1.61555e-07 1.00000e-03 1.61605e-07 1.00000e-03 1.61610e-07 0.00000e+00
+ 1.63550e-07 0.00000e+00 1.63555e-07 1.00000e-03 1.63605e-07 1.00000e-03
+ 1.63610e-07 0.00000e+00 1.65550e-07 0.00000e+00 1.65555e-07 1.00000e-03
+ 1.65605e-07 1.00000e-03 1.65610e-07 0.00000e+00 1.67550e-07 0.00000e+00
+ 1.67555e-07 1.00000e-03 1.67605e-07 1.00000e-03 1.67610e-07 0.00000e+00
+ 1.69550e-07 0.00000e+00 1.69555e-07 1.00000e-03 1.69605e-07 1.00000e-03
+ 1.69610e-07 0.00000e+00 1.71550e-07 0.00000e+00 1.71555e-07 1.00000e-03
+ 1.71605e-07 1.00000e-03 1.71610e-07 0.00000e+00 1.73550e-07 0.00000e+00
+ 1.73555e-07 1.00000e-03 1.73605e-07 1.00000e-03 1.73610e-07 0.00000e+00
+ 1.75550e-07 0.00000e+00 1.75555e-07 1.00000e-03 1.75605e-07 1.00000e-03
+ 1.75610e-07 0.00000e+00 1.77550e-07 0.00000e+00 1.77555e-07 1.00000e-03
+ 1.77605e-07 1.00000e-03 1.77610e-07 0.00000e+00 1.79550e-07 0.00000e+00
+ 1.79555e-07 1.00000e-03 1.79605e-07 1.00000e-03 1.79610e-07 0.00000e+00
+ 1.81550e-07 0.00000e+00 1.81555e-07 1.00000e-03 1.81605e-07 1.00000e-03
+ 1.81610e-07 0.00000e+00 1.83550e-07 0.00000e+00 1.83555e-07 1.00000e-03
+ 1.83605e-07 1.00000e-03 1.83610e-07 0.00000e+00 1.85550e-07 0.00000e+00
+ 1.85555e-07 1.00000e-03 1.85605e-07 1.00000e-03 1.85610e-07 0.00000e+00
+ 1.87550e-07 0.00000e+00 1.87555e-07 1.00000e-03 1.87605e-07 1.00000e-03
+ 1.87610e-07 0.00000e+00 1.89550e-07 0.00000e+00 1.89555e-07 1.00000e-03
+ 1.89605e-07 1.00000e-03 1.89610e-07 0.00000e+00 1.91550e-07 0.00000e+00
+ 1.91555e-07 1.00000e-03 1.91605e-07 1.00000e-03 1.91610e-07 0.00000e+00
+ 1.93550e-07 0.00000e+00 1.93555e-07 1.00000e-03 1.93605e-07 1.00000e-03
+ 1.93610e-07 0.00000e+00 1.95550e-07 0.00000e+00 1.95555e-07 1.00000e-03
+ 1.95605e-07 1.00000e-03 1.95610e-07 0.00000e+00 1.97550e-07 0.00000e+00
+ 1.97555e-07 1.00000e-03 1.97605e-07 1.00000e-03 1.97610e-07 0.00000e+00
+ 1.99550e-07 0.00000e+00 1.99555e-07 1.00000e-03 1.99605e-07 1.00000e-03
+ 1.99610e-07 0.00000e+00)
IIN2 0 IN2 PWL(0 0 20P 0 2.55000e-09 0.00000e+00 2.55500e-09 1.00000e-03 2.60500e-09 1.00000e-03
+ 2.61000e-09 0.00000e+00 3.55000e-09 0.00000e+00 3.55500e-09 1.00000e-03
+ 3.60500e-09 1.00000e-03 3.61000e-09 0.00000e+00 6.55000e-09 0.00000e+00
+ 6.55500e-09 1.00000e-03 6.60500e-09 1.00000e-03 6.61000e-09 0.00000e+00
+ 7.55000e-09 0.00000e+00 7.55500e-09 1.00000e-03 7.60500e-09 1.00000e-03
+ 7.61000e-09 0.00000e+00 1.05500e-08 0.00000e+00 1.05550e-08 1.00000e-03
+ 1.06050e-08 1.00000e-03 1.06100e-08 0.00000e+00 1.15500e-08 0.00000e+00
+ 1.15550e-08 1.00000e-03 1.16050e-08 1.00000e-03 1.16100e-08 0.00000e+00
+ 1.45500e-08 0.00000e+00 1.45550e-08 1.00000e-03 1.46050e-08 1.00000e-03
+ 1.46100e-08 0.00000e+00 1.55500e-08 0.00000e+00 1.55550e-08 1.00000e-03
+ 1.56050e-08 1.00000e-03 1.56100e-08 0.00000e+00 1.85500e-08 0.00000e+00
+ 1.85550e-08 1.00000e-03 1.86050e-08 1.00000e-03 1.86100e-08 0.00000e+00
+ 1.95500e-08 0.00000e+00 1.95550e-08 1.00000e-03 1.96050e-08 1.00000e-03
+ 1.96100e-08 0.00000e+00 2.25500e-08 0.00000e+00 2.25550e-08 1.00000e-03
+ 2.26050e-08 1.00000e-03 2.26100e-08 0.00000e+00 2.35500e-08 0.00000e+00
+ 2.35550e-08 1.00000e-03 2.36050e-08 1.00000e-03 2.36100e-08 0.00000e+00
+ 2.65500e-08 0.00000e+00 2.65550e-08 1.00000e-03 2.66050e-08 1.00000e-03
+ 2.66100e-08 0.00000e+00 2.75500e-08 0.00000e+00 2.75550e-08 1.00000e-03
+ 2.76050e-08 1.00000e-03 2.76100e-08 0.00000e+00 3.05500e-08 0.00000e+00
+ 3.05550e-08 1.00000e-03 3.06050e-08 1.00000e-03 3.06100e-08 0.00000e+00
+ 3.15500e-08 0.00000e+00 3.15550e-08 1.00000e-03 3.16050e-08 1.00000e-03
+ 3.16100e-08 0.00000e+00 3.45500e-08 0.00000e+00 3.45550e-08 1.00000e-03
+ 3.46050e-08 1.00000e-03 3.46100e-08 0.00000e+00 3.55500e-08 0.00000e+00
+ 3.55550e-08 1.00000e-03 3.56050e-08 1.00000e-03 3.56100e-08 0.00000e+00
+ 3.85500e-08 0.00000e+00 3.85550e-08 1.00000e-03 3.86050e-08 1.00000e-03
+ 3.86100e-08 0.00000e+00 3.95500e-08 0.00000e+00 3.95550e-08 1.00000e-03
+ 3.96050e-08 1.00000e-03 3.96100e-08 0.00000e+00 4.25500e-08 0.00000e+00
+ 4.25550e-08 1.00000e-03 4.26050e-08 1.00000e-03 4.26100e-08 0.00000e+00
+ 4.35500e-08 0.00000e+00 4.35550e-08 1.00000e-03 4.36050e-08 1.00000e-03
+ 4.36100e-08 0.00000e+00 4.65500e-08 0.00000e+00 4.65550e-08 1.00000e-03
+ 4.66050e-08 1.00000e-03 4.66100e-08 0.00000e+00 4.75500e-08 0.00000e+00
+ 4.75550e-08 1.00000e-03 4.76050e-08 1.00000e-03 4.76100e-08 0.00000e+00
+ 5.05500e-08 0.00000e+00 5.05550e-08 1.00000e-03 5.06050e-08 1.00000e-03
+ 5.06100e-08 0.00000e+00 5.15500e-08 0.00000e+00 5.15550e-08 1.00000e-03
+ 5.16050e-08 1.00000e-03 5.16100e-08 0.00000e+00 5.45500e-08 0.00000e+00
+ 5.45550e-08 1.00000e-03 5.46050e-08 1.00000e-03 5.46100e-08 0.00000e+00
+ 5.55500e-08 0.00000e+00 5.55550e-08 1.00000e-03 5.56050e-08 1.00000e-03
+ 5.56100e-08 0.00000e+00 5.85500e-08 0.00000e+00 5.85550e-08 1.00000e-03
+ 5.86050e-08 1.00000e-03 5.86100e-08 0.00000e+00 5.95500e-08 0.00000e+00
+ 5.95550e-08 1.00000e-03 5.96050e-08 1.00000e-03 5.96100e-08 0.00000e+00
+ 6.25500e-08 0.00000e+00 6.25550e-08 1.00000e-03 6.26050e-08 1.00000e-03
+ 6.26100e-08 0.00000e+00 6.35500e-08 0.00000e+00 6.35550e-08 1.00000e-03
+ 6.36050e-08 1.00000e-03 6.36100e-08 0.00000e+00 6.65500e-08 0.00000e+00
+ 6.65550e-08 1.00000e-03 6.66050e-08 1.00000e-03 6.66100e-08 0.00000e+00
+ 6.75500e-08 0.00000e+00 6.75550e-08 1.00000e-03 6.76050e-08 1.00000e-03
+ 6.76100e-08 0.00000e+00 7.05500e-08 0.00000e+00 7.05550e-08 1.00000e-03
+ 7.06050e-08 1.00000e-03 7.06100e-08 0.00000e+00 7.15500e-08 0.00000e+00
+ 7.15550e-08 1.00000e-03 7.16050e-08 1.00000e-03 7.16100e-08 0.00000e+00
+ 7.45500e-08 0.00000e+00 7.45550e-08 1.00000e-03 7.46050e-08 1.00000e-03
+ 7.46100e-08 0.00000e+00 7.55500e-08 0.00000e+00 7.55550e-08 1.00000e-03
+ 7.56050e-08 1.00000e-03 7.56100e-08 0.00000e+00 7.85500e-08 0.00000e+00
+ 7.85550e-08 1.00000e-03 7.86050e-08 1.00000e-03 7.86100e-08 0.00000e+00
+ 7.95500e-08 0.00000e+00 7.95550e-08 1.00000e-03 7.96050e-08 1.00000e-03
+ 7.96100e-08 0.00000e+00 8.25500e-08 0.00000e+00 8.25550e-08 1.00000e-03
+ 8.26050e-08 1.00000e-03 8.26100e-08 0.00000e+00 8.35500e-08 0.00000e+00
+ 8.35550e-08 1.00000e-03 8.36050e-08 1.00000e-03 8.36100e-08 0.00000e+00
+ 8.65500e-08 0.00000e+00 8.65550e-08 1.00000e-03 8.66050e-08 1.00000e-03
+ 8.66100e-08 0.00000e+00 8.75500e-08 0.00000e+00 8.75550e-08 1.00000e-03
+ 8.76050e-08 1.00000e-03 8.76100e-08 0.00000e+00 9.05500e-08 0.00000e+00
+ 9.05550e-08 1.00000e-03 9.06050e-08 1.00000e-03 9.06100e-08 0.00000e+00
+ 9.15500e-08 0.00000e+00 9.15550e-08 1.00000e-03 9.16050e-08 1.00000e-03
+ 9.16100e-08 0.00000e+00 9.45500e-08 0.00000e+00 9.45550e-08 1.00000e-03
+ 9.46050e-08 1.00000e-03 9.46100e-08 0.00000e+00 9.55500e-08 0.00000e+00
+ 9.55550e-08 1.00000e-03 9.56050e-08 1.00000e-03 9.56100e-08 0.00000e+00
+ 9.85500e-08 0.00000e+00 9.85550e-08 1.00000e-03 9.86050e-08 1.00000e-03
+ 9.86100e-08 0.00000e+00 9.95500e-08 0.00000e+00 9.95550e-08 1.00000e-03
+ 9.96050e-08 1.00000e-03 9.96100e-08 0.00000e+00 1.02550e-07 0.00000e+00
+ 1.02555e-07 1.00000e-03 1.02605e-07 1.00000e-03 1.02610e-07 0.00000e+00
+ 1.03550e-07 0.00000e+00 1.03555e-07 1.00000e-03 1.03605e-07 1.00000e-03
+ 1.03610e-07 0.00000e+00 1.06550e-07 0.00000e+00 1.06555e-07 1.00000e-03
+ 1.06605e-07 1.00000e-03 1.06610e-07 0.00000e+00 1.07550e-07 0.00000e+00
+ 1.07555e-07 1.00000e-03 1.07605e-07 1.00000e-03 1.07610e-07 0.00000e+00
+ 1.10550e-07 0.00000e+00 1.10555e-07 1.00000e-03 1.10605e-07 1.00000e-03
+ 1.10610e-07 0.00000e+00 1.11550e-07 0.00000e+00 1.11555e-07 1.00000e-03
+ 1.11605e-07 1.00000e-03 1.11610e-07 0.00000e+00 1.14550e-07 0.00000e+00
+ 1.14555e-07 1.00000e-03 1.14605e-07 1.00000e-03 1.14610e-07 0.00000e+00
+ 1.15550e-07 0.00000e+00 1.15555e-07 1.00000e-03 1.15605e-07 1.00000e-03
+ 1.15610e-07 0.00000e+00 1.18550e-07 0.00000e+00 1.18555e-07 1.00000e-03
+ 1.18605e-07 1.00000e-03 1.18610e-07 0.00000e+00 1.19550e-07 0.00000e+00
+ 1.19555e-07 1.00000e-03 1.19605e-07 1.00000e-03 1.19610e-07 0.00000e+00
+ 1.22550e-07 0.00000e+00 1.22555e-07 1.00000e-03 1.22605e-07 1.00000e-03
+ 1.22610e-07 0.00000e+00 1.23550e-07 0.00000e+00 1.23555e-07 1.00000e-03
+ 1.23605e-07 1.00000e-03 1.23610e-07 0.00000e+00 1.26550e-07 0.00000e+00
+ 1.26555e-07 1.00000e-03 1.26605e-07 1.00000e-03 1.26610e-07 0.00000e+00
+ 1.27550e-07 0.00000e+00 1.27555e-07 1.00000e-03 1.27605e-07 1.00000e-03
+ 1.27610e-07 0.00000e+00 1.30550e-07 0.00000e+00 1.30555e-07 1.00000e-03
+ 1.30605e-07 1.00000e-03 1.30610e-07 0.00000e+00 1.31550e-07 0.00000e+00
+ 1.31555e-07 1.00000e-03 1.31605e-07 1.00000e-03 1.31610e-07 0.00000e+00
+ 1.34550e-07 0.00000e+00 1.34555e-07 1.00000e-03 1.34605e-07 1.00000e-03
+ 1.34610e-07 0.00000e+00 1.35550e-07 0.00000e+00 1.35555e-07 1.00000e-03
+ 1.35605e-07 1.00000e-03 1.35610e-07 0.00000e+00 1.38550e-07 0.00000e+00
+ 1.38555e-07 1.00000e-03 1.38605e-07 1.00000e-03 1.38610e-07 0.00000e+00
+ 1.39550e-07 0.00000e+00 1.39555e-07 1.00000e-03 1.39605e-07 1.00000e-03
+ 1.39610e-07 0.00000e+00 1.42550e-07 0.00000e+00 1.42555e-07 1.00000e-03
+ 1.42605e-07 1.00000e-03 1.42610e-07 0.00000e+00 1.43550e-07 0.00000e+00
+ 1.43555e-07 1.00000e-03 1.43605e-07 1.00000e-03 1.43610e-07 0.00000e+00
+ 1.46550e-07 0.00000e+00 1.46555e-07 1.00000e-03 1.46605e-07 1.00000e-03
+ 1.46610e-07 0.00000e+00 1.47550e-07 0.00000e+00 1.47555e-07 1.00000e-03
+ 1.47605e-07 1.00000e-03 1.47610e-07 0.00000e+00 1.50550e-07 0.00000e+00
+ 1.50555e-07 1.00000e-03 1.50605e-07 1.00000e-03 1.50610e-07 0.00000e+00
+ 1.51550e-07 0.00000e+00 1.51555e-07 1.00000e-03 1.51605e-07 1.00000e-03
+ 1.51610e-07 0.00000e+00 1.54550e-07 0.00000e+00 1.54555e-07 1.00000e-03
+ 1.54605e-07 1.00000e-03 1.54610e-07 0.00000e+00 1.55550e-07 0.00000e+00
+ 1.55555e-07 1.00000e-03 1.55605e-07 1.00000e-03 1.55610e-07 0.00000e+00
+ 1.58550e-07 0.00000e+00 1.58555e-07 1.00000e-03 1.58605e-07 1.00000e-03
+ 1.58610e-07 0.00000e+00 1.59550e-07 0.00000e+00 1.59555e-07 1.00000e-03
+ 1.59605e-07 1.00000e-03 1.59610e-07 0.00000e+00 1.62550e-07 0.00000e+00
+ 1.62555e-07 1.00000e-03 1.62605e-07 1.00000e-03 1.62610e-07 0.00000e+00
+ 1.63550e-07 0.00000e+00 1.63555e-07 1.00000e-03 1.63605e-07 1.00000e-03
+ 1.63610e-07 0.00000e+00 1.66550e-07 0.00000e+00 1.66555e-07 1.00000e-03
+ 1.66605e-07 1.00000e-03 1.66610e-07 0.00000e+00 1.67550e-07 0.00000e+00
+ 1.67555e-07 1.00000e-03 1.67605e-07 1.00000e-03 1.67610e-07 0.00000e+00
+ 1.70550e-07 0.00000e+00 1.70555e-07 1.00000e-03 1.70605e-07 1.00000e-03
+ 1.70610e-07 0.00000e+00 1.71550e-07 0.00000e+00 1.71555e-07 1.00000e-03
+ 1.71605e-07 1.00000e-03 1.71610e-07 0.00000e+00 1.74550e-07 0.00000e+00
+ 1.74555e-07 1.00000e-03 1.74605e-07 1.00000e-03 1.74610e-07 0.00000e+00
+ 1.75550e-07 0.00000e+00 1.75555e-07 1.00000e-03 1.75605e-07 1.00000e-03
+ 1.75610e-07 0.00000e+00 1.78550e-07 0.00000e+00 1.78555e-07 1.00000e-03
+ 1.78605e-07 1.00000e-03 1.78610e-07 0.00000e+00 1.79550e-07 0.00000e+00
+ 1.79555e-07 1.00000e-03 1.79605e-07 1.00000e-03 1.79610e-07 0.00000e+00
+ 1.82550e-07 0.00000e+00 1.82555e-07 1.00000e-03 1.82605e-07 1.00000e-03
+ 1.82610e-07 0.00000e+00 1.83550e-07 0.00000e+00 1.83555e-07 1.00000e-03
+ 1.83605e-07 1.00000e-03 1.83610e-07 0.00000e+00 1.86550e-07 0.00000e+00
+ 1.86555e-07 1.00000e-03 1.86605e-07 1.00000e-03 1.86610e-07 0.00000e+00
+ 1.87550e-07 0.00000e+00 1.87555e-07 1.00000e-03 1.87605e-07 1.00000e-03
+ 1.87610e-07 0.00000e+00 1.90550e-07 0.00000e+00 1.90555e-07 1.00000e-03
+ 1.90605e-07 1.00000e-03 1.90610e-07 0.00000e+00 1.91550e-07 0.00000e+00
+ 1.91555e-07 1.00000e-03 1.91605e-07 1.00000e-03 1.91610e-07 0.00000e+00
+ 1.94550e-07 0.00000e+00 1.94555e-07 1.00000e-03 1.94605e-07 1.00000e-03
+ 1.94610e-07 0.00000e+00 1.95550e-07 0.00000e+00 1.95555e-07 1.00000e-03
+ 1.95605e-07 1.00000e-03 1.95610e-07 0.00000e+00 1.98550e-07 0.00000e+00
+ 1.98555e-07 1.00000e-03 1.98605e-07 1.00000e-03 1.98610e-07 0.00000e+00
+ 1.99550e-07 0.00000e+00 1.99555e-07 1.00000e-03 1.99605e-07 1.00000e-03
+ 1.99610e-07 0.00000e+00)
IINBIAS1 0 INB11 pulse(0 0.001 550p 5p 5p 50p 1000p)
ITARGET 0 TARGET0  PWL(0 0 20P 0 5.50000e-10 0.00000e+00 5.55000e-10 1.00000e-03 6.05000e-10 1.00000e-03
+ 6.10000e-10 0.00000e+00 3.55000e-09 0.00000e+00 3.55500e-09 1.00000e-03
+ 3.60500e-09 1.00000e-03 3.61000e-09 0.00000e+00 4.55000e-09 0.00000e+00
+ 4.55500e-09 1.00000e-03 4.60500e-09 1.00000e-03 4.61000e-09 0.00000e+00
+ 7.55000e-09 0.00000e+00 7.55500e-09 1.00000e-03 7.60500e-09 1.00000e-03
+ 7.61000e-09 0.00000e+00 8.55000e-09 0.00000e+00 8.55500e-09 1.00000e-03
+ 8.60500e-09 1.00000e-03 8.61000e-09 0.00000e+00 1.15500e-08 0.00000e+00
+ 1.15550e-08 1.00000e-03 1.16050e-08 1.00000e-03 1.16100e-08 0.00000e+00
+ 1.25500e-08 0.00000e+00 1.25550e-08 1.00000e-03 1.26050e-08 1.00000e-03
+ 1.26100e-08 0.00000e+00 1.55500e-08 0.00000e+00 1.55550e-08 1.00000e-03
+ 1.56050e-08 1.00000e-03 1.56100e-08 0.00000e+00 1.65500e-08 0.00000e+00
+ 1.65550e-08 1.00000e-03 1.66050e-08 1.00000e-03 1.66100e-08 0.00000e+00
+ 1.95500e-08 0.00000e+00 1.95550e-08 1.00000e-03 1.96050e-08 1.00000e-03
+ 1.96100e-08 0.00000e+00 2.05500e-08 0.00000e+00 2.05550e-08 1.00000e-03
+ 2.06050e-08 1.00000e-03 2.06100e-08 0.00000e+00 2.35500e-08 0.00000e+00
+ 2.35550e-08 1.00000e-03 2.36050e-08 1.00000e-03 2.36100e-08 0.00000e+00
+ 2.45500e-08 0.00000e+00 2.45550e-08 1.00000e-03 2.46050e-08 1.00000e-03
+ 2.46100e-08 0.00000e+00 2.75500e-08 0.00000e+00 2.75550e-08 1.00000e-03
+ 2.76050e-08 1.00000e-03 2.76100e-08 0.00000e+00 2.85500e-08 0.00000e+00
+ 2.85550e-08 1.00000e-03 2.86050e-08 1.00000e-03 2.86100e-08 0.00000e+00
+ 3.15500e-08 0.00000e+00 3.15550e-08 1.00000e-03 3.16050e-08 1.00000e-03
+ 3.16100e-08 0.00000e+00 3.25500e-08 0.00000e+00 3.25550e-08 1.00000e-03
+ 3.26050e-08 1.00000e-03 3.26100e-08 0.00000e+00 3.55500e-08 0.00000e+00
+ 3.55550e-08 1.00000e-03 3.56050e-08 1.00000e-03 3.56100e-08 0.00000e+00
+ 3.65500e-08 0.00000e+00 3.65550e-08 1.00000e-03 3.66050e-08 1.00000e-03
+ 3.66100e-08 0.00000e+00 3.95500e-08 0.00000e+00 3.95550e-08 1.00000e-03
+ 3.96050e-08 1.00000e-03 3.96100e-08 0.00000e+00 4.05500e-08 0.00000e+00
+ 4.05550e-08 1.00000e-03 4.06050e-08 1.00000e-03 4.06100e-08 0.00000e+00
+ 4.35500e-08 0.00000e+00 4.35550e-08 1.00000e-03 4.36050e-08 1.00000e-03
+ 4.36100e-08 0.00000e+00 4.45500e-08 0.00000e+00 4.45550e-08 1.00000e-03
+ 4.46050e-08 1.00000e-03 4.46100e-08 0.00000e+00 4.75500e-08 0.00000e+00
+ 4.75550e-08 1.00000e-03 4.76050e-08 1.00000e-03 4.76100e-08 0.00000e+00
+ 4.85500e-08 0.00000e+00 4.85550e-08 1.00000e-03 4.86050e-08 1.00000e-03
+ 4.86100e-08 0.00000e+00 5.15500e-08 0.00000e+00 5.15550e-08 1.00000e-03
+ 5.16050e-08 1.00000e-03 5.16100e-08 0.00000e+00 5.25500e-08 0.00000e+00
+ 5.25550e-08 1.00000e-03 5.26050e-08 1.00000e-03 5.26100e-08 0.00000e+00
+ 5.55500e-08 0.00000e+00 5.55550e-08 1.00000e-03 5.56050e-08 1.00000e-03
+ 5.56100e-08 0.00000e+00 5.65500e-08 0.00000e+00 5.65550e-08 1.00000e-03
+ 5.66050e-08 1.00000e-03 5.66100e-08 0.00000e+00 5.95500e-08 0.00000e+00
+ 5.95550e-08 1.00000e-03 5.96050e-08 1.00000e-03 5.96100e-08 0.00000e+00
+ 6.05500e-08 0.00000e+00 6.05550e-08 1.00000e-03 6.06050e-08 1.00000e-03
+ 6.06100e-08 0.00000e+00 6.35500e-08 0.00000e+00 6.35550e-08 1.00000e-03
+ 6.36050e-08 1.00000e-03 6.36100e-08 0.00000e+00 6.45500e-08 0.00000e+00
+ 6.45550e-08 1.00000e-03 6.46050e-08 1.00000e-03 6.46100e-08 0.00000e+00
+ 6.75500e-08 0.00000e+00 6.75550e-08 1.00000e-03 6.76050e-08 1.00000e-03
+ 6.76100e-08 0.00000e+00 6.85500e-08 0.00000e+00 6.85550e-08 1.00000e-03
+ 6.86050e-08 1.00000e-03 6.86100e-08 0.00000e+00 7.15500e-08 0.00000e+00
+ 7.15550e-08 1.00000e-03 7.16050e-08 1.00000e-03 7.16100e-08 0.00000e+00
+ 7.25500e-08 0.00000e+00 7.25550e-08 1.00000e-03 7.26050e-08 1.00000e-03
+ 7.26100e-08 0.00000e+00 7.55500e-08 0.00000e+00 7.55550e-08 1.00000e-03
+ 7.56050e-08 1.00000e-03 7.56100e-08 0.00000e+00 7.65500e-08 0.00000e+00
+ 7.65550e-08 1.00000e-03 7.66050e-08 1.00000e-03 7.66100e-08 0.00000e+00
+ 7.95500e-08 0.00000e+00 7.95550e-08 1.00000e-03 7.96050e-08 1.00000e-03
+ 7.96100e-08 0.00000e+00 8.05500e-08 0.00000e+00 8.05550e-08 1.00000e-03
+ 8.06050e-08 1.00000e-03 8.06100e-08 0.00000e+00 8.35500e-08 0.00000e+00
+ 8.35550e-08 1.00000e-03 8.36050e-08 1.00000e-03 8.36100e-08 0.00000e+00
+ 8.45500e-08 0.00000e+00 8.45550e-08 1.00000e-03 8.46050e-08 1.00000e-03
+ 8.46100e-08 0.00000e+00 8.75500e-08 0.00000e+00 8.75550e-08 1.00000e-03
+ 8.76050e-08 1.00000e-03 8.76100e-08 0.00000e+00 8.85500e-08 0.00000e+00
+ 8.85550e-08 1.00000e-03 8.86050e-08 1.00000e-03 8.86100e-08 0.00000e+00
+ 9.15500e-08 0.00000e+00 9.15550e-08 1.00000e-03 9.16050e-08 1.00000e-03
+ 9.16100e-08 0.00000e+00 9.25500e-08 0.00000e+00 9.25550e-08 1.00000e-03
+ 9.26050e-08 1.00000e-03 9.26100e-08 0.00000e+00 9.55500e-08 0.00000e+00
+ 9.55550e-08 1.00000e-03 9.56050e-08 1.00000e-03 9.56100e-08 0.00000e+00
+ 9.65500e-08 0.00000e+00 9.65550e-08 1.00000e-03 9.66050e-08 1.00000e-03
+ 9.66100e-08 0.00000e+00 9.95500e-08 0.00000e+00 9.95550e-08 1.00000e-03
+ 9.96050e-08 1.00000e-03 9.96100e-08 0.00000e+00 1.00550e-07 0.00000e+00
+ 1.00555e-07 1.00000e-03 1.00605e-07 1.00000e-03 1.00610e-07 0.00000e+00
+ 1.03550e-07 0.00000e+00 1.03555e-07 1.00000e-03 1.03605e-07 1.00000e-03
+ 1.03610e-07 0.00000e+00 1.04550e-07 0.00000e+00 1.04555e-07 1.00000e-03
+ 1.04605e-07 1.00000e-03 1.04610e-07 0.00000e+00 1.07550e-07 0.00000e+00
+ 1.07555e-07 1.00000e-03 1.07605e-07 1.00000e-03 1.07610e-07 0.00000e+00
+ 1.08550e-07 0.00000e+00 1.08555e-07 1.00000e-03 1.08605e-07 1.00000e-03
+ 1.08610e-07 0.00000e+00 1.11550e-07 0.00000e+00 1.11555e-07 1.00000e-03
+ 1.11605e-07 1.00000e-03 1.11610e-07 0.00000e+00 1.12550e-07 0.00000e+00
+ 1.12555e-07 1.00000e-03 1.12605e-07 1.00000e-03 1.12610e-07 0.00000e+00
+ 1.15550e-07 0.00000e+00 1.15555e-07 1.00000e-03 1.15605e-07 1.00000e-03
+ 1.15610e-07 0.00000e+00 1.16550e-07 0.00000e+00 1.16555e-07 1.00000e-03
+ 1.16605e-07 1.00000e-03 1.16610e-07 0.00000e+00 1.19550e-07 0.00000e+00
+ 1.19555e-07 1.00000e-03 1.19605e-07 1.00000e-03 1.19610e-07 0.00000e+00
+ 1.20550e-07 0.00000e+00 1.20555e-07 1.00000e-03 1.20605e-07 1.00000e-03
+ 1.20610e-07 0.00000e+00 1.23550e-07 0.00000e+00 1.23555e-07 1.00000e-03
+ 1.23605e-07 1.00000e-03 1.23610e-07 0.00000e+00 1.24550e-07 0.00000e+00
+ 1.24555e-07 1.00000e-03 1.24605e-07 1.00000e-03 1.24610e-07 0.00000e+00
+ 1.27550e-07 0.00000e+00 1.27555e-07 1.00000e-03 1.27605e-07 1.00000e-03
+ 1.27610e-07 0.00000e+00 1.28550e-07 0.00000e+00 1.28555e-07 1.00000e-03
+ 1.28605e-07 1.00000e-03 1.28610e-07 0.00000e+00 1.31550e-07 0.00000e+00
+ 1.31555e-07 1.00000e-03 1.31605e-07 1.00000e-03 1.31610e-07 0.00000e+00
+ 1.32550e-07 0.00000e+00 1.32555e-07 1.00000e-03 1.32605e-07 1.00000e-03
+ 1.32610e-07 0.00000e+00 1.35550e-07 0.00000e+00 1.35555e-07 1.00000e-03
+ 1.35605e-07 1.00000e-03 1.35610e-07 0.00000e+00 1.36550e-07 0.00000e+00
+ 1.36555e-07 1.00000e-03 1.36605e-07 1.00000e-03 1.36610e-07 0.00000e+00
+ 1.39550e-07 0.00000e+00 1.39555e-07 1.00000e-03 1.39605e-07 1.00000e-03
+ 1.39610e-07 0.00000e+00 1.40550e-07 0.00000e+00 1.40555e-07 1.00000e-03
+ 1.40605e-07 1.00000e-03 1.40610e-07 0.00000e+00 1.43550e-07 0.00000e+00
+ 1.43555e-07 1.00000e-03 1.43605e-07 1.00000e-03 1.43610e-07 0.00000e+00
+ 1.44550e-07 0.00000e+00 1.44555e-07 1.00000e-03 1.44605e-07 1.00000e-03
+ 1.44610e-07 0.00000e+00 1.47550e-07 0.00000e+00 1.47555e-07 1.00000e-03
+ 1.47605e-07 1.00000e-03 1.47610e-07 0.00000e+00 1.48550e-07 0.00000e+00
+ 1.48555e-07 1.00000e-03 1.48605e-07 1.00000e-03 1.48610e-07 0.00000e+00
+ 1.51550e-07 0.00000e+00 1.51555e-07 1.00000e-03 1.51605e-07 1.00000e-03
+ 1.51610e-07 0.00000e+00 1.52550e-07 0.00000e+00 1.52555e-07 1.00000e-03
+ 1.52605e-07 1.00000e-03 1.52610e-07 0.00000e+00 1.55550e-07 0.00000e+00
+ 1.55555e-07 1.00000e-03 1.55605e-07 1.00000e-03 1.55610e-07 0.00000e+00
+ 1.56550e-07 0.00000e+00 1.56555e-07 1.00000e-03 1.56605e-07 1.00000e-03
+ 1.56610e-07 0.00000e+00 1.59550e-07 0.00000e+00 1.59555e-07 1.00000e-03
+ 1.59605e-07 1.00000e-03 1.59610e-07 0.00000e+00 1.60550e-07 0.00000e+00
+ 1.60555e-07 1.00000e-03 1.60605e-07 1.00000e-03 1.60610e-07 0.00000e+00
+ 1.63550e-07 0.00000e+00 1.63555e-07 1.00000e-03 1.63605e-07 1.00000e-03
+ 1.63610e-07 0.00000e+00 1.64550e-07 0.00000e+00 1.64555e-07 1.00000e-03
+ 1.64605e-07 1.00000e-03 1.64610e-07 0.00000e+00 1.67550e-07 0.00000e+00
+ 1.67555e-07 1.00000e-03 1.67605e-07 1.00000e-03 1.67610e-07 0.00000e+00
+ 1.68550e-07 0.00000e+00 1.68555e-07 1.00000e-03 1.68605e-07 1.00000e-03
+ 1.68610e-07 0.00000e+00 1.71550e-07 0.00000e+00 1.71555e-07 1.00000e-03
+ 1.71605e-07 1.00000e-03 1.71610e-07 0.00000e+00 1.72550e-07 0.00000e+00
+ 1.72555e-07 1.00000e-03 1.72605e-07 1.00000e-03 1.72610e-07 0.00000e+00
+ 1.75550e-07 0.00000e+00 1.75555e-07 1.00000e-03 1.75605e-07 1.00000e-03
+ 1.75610e-07 0.00000e+00 1.76550e-07 0.00000e+00 1.76555e-07 1.00000e-03
+ 1.76605e-07 1.00000e-03 1.76610e-07 0.00000e+00 1.79550e-07 0.00000e+00
+ 1.79555e-07 1.00000e-03 1.79605e-07 1.00000e-03 1.79610e-07 0.00000e+00
+ 1.80550e-07 0.00000e+00 1.80555e-07 1.00000e-03 1.80605e-07 1.00000e-03
+ 1.80610e-07 0.00000e+00 1.83550e-07 0.00000e+00 1.83555e-07 1.00000e-03
+ 1.83605e-07 1.00000e-03 1.83610e-07 0.00000e+00 1.84550e-07 0.00000e+00
+ 1.84555e-07 1.00000e-03 1.84605e-07 1.00000e-03 1.84610e-07 0.00000e+00
+ 1.87550e-07 0.00000e+00 1.87555e-07 1.00000e-03 1.87605e-07 1.00000e-03
+ 1.87610e-07 0.00000e+00 1.88550e-07 0.00000e+00 1.88555e-07 1.00000e-03
+ 1.88605e-07 1.00000e-03 1.88610e-07 0.00000e+00 1.91550e-07 0.00000e+00
+ 1.91555e-07 1.00000e-03 1.91605e-07 1.00000e-03 1.91610e-07 0.00000e+00
+ 1.92550e-07 0.00000e+00 1.92555e-07 1.00000e-03 1.92605e-07 1.00000e-03
+ 1.92610e-07 0.00000e+00 1.95550e-07 0.00000e+00 1.95555e-07 1.00000e-03
+ 1.95605e-07 1.00000e-03 1.95610e-07 0.00000e+00 1.96550e-07 0.00000e+00
+ 1.96555e-07 1.00000e-03 1.96605e-07 1.00000e-03 1.96610e-07 0.00000e+00
+ 1.99550e-07 0.00000e+00 1.99555e-07 1.00000e-03 1.99605e-07 1.00000e-03
+ 1.99610e-07 0.00000e+00)
Iactualsynbias21 0 ACTUALSYNB21x PWL(0 0 6.40000e-10 0.00000e+00 6.65000e-10 6.70000e-04 7.00000e-10 0.00000e+00
+ 8.40000e-10 0.00000e+00 8.65000e-10 6.70000e-04 9.00000e-10 0.00000e+00
+ 1.04000e-09 0.00000e+00 1.06500e-09 6.70000e-04 1.10000e-09 0.00000e+00
+ 1.24000e-09 0.00000e+00 1.26500e-09 6.70000e-04 1.30000e-09 0.00000e+00
+ 1.44000e-09 0.00000e+00 1.46500e-09 6.70000e-04 1.50000e-09 0.00000e+00
+ 1.64000e-09 0.00000e+00 1.66500e-09 6.70000e-04 1.70000e-09 0.00000e+00
+ 1.84000e-09 0.00000e+00 1.86500e-09 6.70000e-04 1.90000e-09 0.00000e+00
+ 2.04000e-09 0.00000e+00 2.06500e-09 6.70000e-04 2.10000e-09 0.00000e+00
+ 2.24000e-09 0.00000e+00 2.26500e-09 6.70000e-04 2.30000e-09 0.00000e+00
+ 2.44000e-09 0.00000e+00 2.46500e-09 6.70000e-04 2.50000e-09 0.00000e+00
+ 2.64000e-09 0.00000e+00 2.66500e-09 6.70000e-04 2.70000e-09 0.00000e+00
+ 2.84000e-09 0.00000e+00 2.86500e-09 6.70000e-04 2.90000e-09 0.00000e+00
+ 3.04000e-09 0.00000e+00 3.06500e-09 6.70000e-04 3.10000e-09 0.00000e+00
+ 3.24000e-09 0.00000e+00 3.26500e-09 6.70000e-04 3.30000e-09 0.00000e+00
+ 3.44000e-09 0.00000e+00 3.46500e-09 6.70000e-04 3.50000e-09 0.00000e+00
+ 3.64000e-09 0.00000e+00 3.66500e-09 6.70000e-04 3.70000e-09 0.00000e+00
+ 3.84000e-09 0.00000e+00 3.86500e-09 6.70000e-04 3.90000e-09 0.00000e+00
+ 4.04000e-09 0.00000e+00 4.06500e-09 6.70000e-04 4.10000e-09 0.00000e+00
+ 4.24000e-09 0.00000e+00 4.26500e-09 6.70000e-04 4.30000e-09 0.00000e+00
+ 4.44000e-09 0.00000e+00 4.46500e-09 6.70000e-04 4.50000e-09 0.00000e+00
+ 4.64000e-09 0.00000e+00 4.66500e-09 6.70000e-04 4.70000e-09 0.00000e+00
+ 4.84000e-09 0.00000e+00 4.86500e-09 6.70000e-04 4.90000e-09 0.00000e+00
+ 5.04000e-09 0.00000e+00 5.06500e-09 6.70000e-04 5.10000e-09 0.00000e+00
+ 5.24000e-09 0.00000e+00 5.26500e-09 6.70000e-04 5.30000e-09 0.00000e+00
+ 5.44000e-09 0.00000e+00 5.46500e-09 6.70000e-04 5.50000e-09 0.00000e+00
+ 5.64000e-09 0.00000e+00 5.66500e-09 6.70000e-04 5.70000e-09 0.00000e+00
+ 5.84000e-09 0.00000e+00 5.86500e-09 6.70000e-04 5.90000e-09 0.00000e+00
+ 6.04000e-09 0.00000e+00 6.06500e-09 6.70000e-04 6.10000e-09 0.00000e+00
+ 6.24000e-09 0.00000e+00 6.26500e-09 6.70000e-04 6.30000e-09 0.00000e+00
+ 6.44000e-09 0.00000e+00 6.46500e-09 6.70000e-04 6.50000e-09 0.00000e+00
+ 6.64000e-09 0.00000e+00 6.66500e-09 6.70000e-04 6.70000e-09 0.00000e+00
+ 6.84000e-09 0.00000e+00 6.86500e-09 6.70000e-04 6.90000e-09 0.00000e+00
+ 7.04000e-09 0.00000e+00 7.06500e-09 6.70000e-04 7.10000e-09 0.00000e+00
+ 7.24000e-09 0.00000e+00 7.26500e-09 6.70000e-04 7.30000e-09 0.00000e+00
+ 7.44000e-09 0.00000e+00 7.46500e-09 6.70000e-04 7.50000e-09 0.00000e+00
+ 7.64000e-09 0.00000e+00 7.66500e-09 6.70000e-04 7.70000e-09 0.00000e+00
+ 7.84000e-09 0.00000e+00 7.86500e-09 6.70000e-04 7.90000e-09 0.00000e+00
+ 8.04000e-09 0.00000e+00 8.06500e-09 6.70000e-04 8.10000e-09 0.00000e+00
+ 8.24000e-09 0.00000e+00 8.26500e-09 6.70000e-04 8.30000e-09 0.00000e+00
+ 8.44000e-09 0.00000e+00 8.46500e-09 6.70000e-04 8.50000e-09 0.00000e+00
+ 8.64000e-09 0.00000e+00 8.66500e-09 6.70000e-04 8.70000e-09 0.00000e+00
+ 8.84000e-09 0.00000e+00 8.86500e-09 6.70000e-04 8.90000e-09 0.00000e+00
+ 9.04000e-09 0.00000e+00 9.06500e-09 6.70000e-04 9.10000e-09 0.00000e+00
+ 9.24000e-09 0.00000e+00 9.26500e-09 6.70000e-04 9.30000e-09 0.00000e+00
+ 9.44000e-09 0.00000e+00 9.46500e-09 6.70000e-04 9.50000e-09 0.00000e+00
+ 9.64000e-09 0.00000e+00 9.66500e-09 6.70000e-04 9.70000e-09 0.00000e+00
+ 9.84000e-09 0.00000e+00 9.86500e-09 6.70000e-04 9.90000e-09 0.00000e+00
+ 1.00400e-08 0.00000e+00 1.00650e-08 6.70000e-04 1.01000e-08 0.00000e+00
+ 1.02400e-08 0.00000e+00 1.02650e-08 6.70000e-04 1.03000e-08 0.00000e+00
+ 1.04400e-08 0.00000e+00 1.04650e-08 6.70000e-04 1.05000e-08 0.00000e+00
+ 1.06400e-08 0.00000e+00 1.06650e-08 6.70000e-04 1.07000e-08 0.00000e+00
+ 1.08400e-08 0.00000e+00 1.08650e-08 6.70000e-04 1.09000e-08 0.00000e+00
+ 1.10400e-08 0.00000e+00 1.10650e-08 6.70000e-04 1.11000e-08 0.00000e+00
+ 1.12400e-08 0.00000e+00 1.12650e-08 6.70000e-04 1.13000e-08 0.00000e+00
+ 1.14400e-08 0.00000e+00 1.14650e-08 6.70000e-04 1.15000e-08 0.00000e+00
+ 1.16400e-08 0.00000e+00 1.16650e-08 6.70000e-04 1.17000e-08 0.00000e+00
+ 1.18400e-08 0.00000e+00 1.18650e-08 6.70000e-04 1.19000e-08 0.00000e+00
+ 1.20400e-08 0.00000e+00 1.20650e-08 6.70000e-04 1.21000e-08 0.00000e+00
+ 1.22400e-08 0.00000e+00 1.22650e-08 6.70000e-04 1.23000e-08 0.00000e+00
+ 1.24400e-08 0.00000e+00 1.24650e-08 6.70000e-04 1.25000e-08 0.00000e+00
+ 1.26400e-08 0.00000e+00 1.26650e-08 6.70000e-04 1.27000e-08 0.00000e+00
+ 1.28400e-08 0.00000e+00 1.28650e-08 6.70000e-04 1.29000e-08 0.00000e+00
+ 1.30400e-08 0.00000e+00 1.30650e-08 6.70000e-04 1.31000e-08 0.00000e+00
+ 1.32400e-08 0.00000e+00 1.32650e-08 6.70000e-04 1.33000e-08 0.00000e+00
+ 1.34400e-08 0.00000e+00 1.34650e-08 6.70000e-04 1.35000e-08 0.00000e+00
+ 1.36400e-08 0.00000e+00 1.36650e-08 6.70000e-04 1.37000e-08 0.00000e+00
+ 1.38400e-08 0.00000e+00 1.38650e-08 6.70000e-04 1.39000e-08 0.00000e+00
+ 1.40400e-08 0.00000e+00 1.40650e-08 6.70000e-04 1.41000e-08 0.00000e+00
+ 1.42400e-08 0.00000e+00 1.42650e-08 6.70000e-04 1.43000e-08 0.00000e+00
+ 1.44400e-08 0.00000e+00 1.44650e-08 6.70000e-04 1.45000e-08 0.00000e+00
+ 1.46400e-08 0.00000e+00 1.46650e-08 6.70000e-04 1.47000e-08 0.00000e+00
+ 1.48400e-08 0.00000e+00 1.48650e-08 6.70000e-04 1.49000e-08 0.00000e+00
+ 1.50400e-08 0.00000e+00 1.50650e-08 6.70000e-04 1.51000e-08 0.00000e+00
+ 1.52400e-08 0.00000e+00 1.52650e-08 6.70000e-04 1.53000e-08 0.00000e+00
+ 1.54400e-08 0.00000e+00 1.54650e-08 6.70000e-04 1.55000e-08 0.00000e+00
+ 1.56400e-08 0.00000e+00 1.56650e-08 6.70000e-04 1.57000e-08 0.00000e+00
+ 1.58400e-08 0.00000e+00 1.58650e-08 6.70000e-04 1.59000e-08 0.00000e+00
+ 1.60400e-08 0.00000e+00 1.60650e-08 6.70000e-04 1.61000e-08 0.00000e+00
+ 1.62400e-08 0.00000e+00 1.62650e-08 6.70000e-04 1.63000e-08 0.00000e+00
+ 1.64400e-08 0.00000e+00 1.64650e-08 6.70000e-04 1.65000e-08 0.00000e+00
+ 1.66400e-08 0.00000e+00 1.66650e-08 6.70000e-04 1.67000e-08 0.00000e+00
+ 1.68400e-08 0.00000e+00 1.68650e-08 6.70000e-04 1.69000e-08 0.00000e+00
+ 1.70400e-08 0.00000e+00 1.70650e-08 6.70000e-04 1.71000e-08 0.00000e+00
+ 1.72400e-08 0.00000e+00 1.72650e-08 6.70000e-04 1.73000e-08 0.00000e+00
+ 1.74400e-08 0.00000e+00 1.74650e-08 6.70000e-04 1.75000e-08 0.00000e+00
+ 1.76400e-08 0.00000e+00 1.76650e-08 6.70000e-04 1.77000e-08 0.00000e+00
+ 1.78400e-08 0.00000e+00 1.78650e-08 6.70000e-04 1.79000e-08 0.00000e+00
+ 1.80400e-08 0.00000e+00 1.80650e-08 6.70000e-04 1.81000e-08 0.00000e+00
+ 1.82400e-08 0.00000e+00 1.82650e-08 6.70000e-04 1.83000e-08 0.00000e+00
+ 1.84400e-08 0.00000e+00 1.84650e-08 6.70000e-04 1.85000e-08 0.00000e+00
+ 1.86400e-08 0.00000e+00 1.86650e-08 6.70000e-04 1.87000e-08 0.00000e+00
+ 1.88400e-08 0.00000e+00 1.88650e-08 6.70000e-04 1.89000e-08 0.00000e+00
+ 1.90400e-08 0.00000e+00 1.90650e-08 6.70000e-04 1.91000e-08 0.00000e+00
+ 1.92400e-08 0.00000e+00 1.92650e-08 6.70000e-04 1.93000e-08 0.00000e+00
+ 1.94400e-08 0.00000e+00 1.94650e-08 6.70000e-04 1.95000e-08 0.00000e+00
+ 1.96400e-08 0.00000e+00 1.96650e-08 6.70000e-04 1.97000e-08 0.00000e+00
+ 1.98400e-08 0.00000e+00 1.98650e-08 6.70000e-04 1.99000e-08 0.00000e+00
+ 2.00400e-08 0.00000e+00 2.00650e-08 6.70000e-04 2.01000e-08 0.00000e+00
+ 2.02400e-08 0.00000e+00 2.02650e-08 6.70000e-04 2.03000e-08 0.00000e+00
+ 2.04400e-08 0.00000e+00 2.04650e-08 6.70000e-04 2.05000e-08 0.00000e+00
+ 2.06400e-08 0.00000e+00 2.06650e-08 6.70000e-04 2.07000e-08 0.00000e+00
+ 2.08400e-08 0.00000e+00 2.08650e-08 6.70000e-04 2.09000e-08 0.00000e+00
+ 2.10400e-08 0.00000e+00 2.10650e-08 6.70000e-04 2.11000e-08 0.00000e+00
+ 2.12400e-08 0.00000e+00 2.12650e-08 6.70000e-04 2.13000e-08 0.00000e+00
+ 2.14400e-08 0.00000e+00 2.14650e-08 6.70000e-04 2.15000e-08 0.00000e+00
+ 2.16400e-08 0.00000e+00 2.16650e-08 6.70000e-04 2.17000e-08 0.00000e+00
+ 2.18400e-08 0.00000e+00 2.18650e-08 6.70000e-04 2.19000e-08 0.00000e+00
+ 2.20400e-08 0.00000e+00 2.20650e-08 6.70000e-04 2.21000e-08 0.00000e+00
+ 2.22400e-08 0.00000e+00 2.22650e-08 6.70000e-04 2.23000e-08 0.00000e+00
+ 2.24400e-08 0.00000e+00 2.24650e-08 6.70000e-04 2.25000e-08 0.00000e+00
+ 2.26400e-08 0.00000e+00 2.26650e-08 6.70000e-04 2.27000e-08 0.00000e+00
+ 2.28400e-08 0.00000e+00 2.28650e-08 6.70000e-04 2.29000e-08 0.00000e+00
+ 2.30400e-08 0.00000e+00 2.30650e-08 6.70000e-04 2.31000e-08 0.00000e+00
+ 2.32400e-08 0.00000e+00 2.32650e-08 6.70000e-04 2.33000e-08 0.00000e+00
+ 2.34400e-08 0.00000e+00 2.34650e-08 6.70000e-04 2.35000e-08 0.00000e+00
+ 2.36400e-08 0.00000e+00 2.36650e-08 6.70000e-04 2.37000e-08 0.00000e+00
+ 2.38400e-08 0.00000e+00 2.38650e-08 6.70000e-04 2.39000e-08 0.00000e+00
+ 2.40400e-08 0.00000e+00 2.40650e-08 6.70000e-04 2.41000e-08 0.00000e+00
+ 2.42400e-08 0.00000e+00 2.42650e-08 6.70000e-04 2.43000e-08 0.00000e+00
+ 2.44400e-08 0.00000e+00 2.44650e-08 6.70000e-04 2.45000e-08 0.00000e+00
+ 2.46400e-08 0.00000e+00 2.46650e-08 6.70000e-04 2.47000e-08 0.00000e+00
+ 2.48400e-08 0.00000e+00 2.48650e-08 6.70000e-04 2.49000e-08 0.00000e+00
+ 2.50400e-08 0.00000e+00 2.50650e-08 6.70000e-04 2.51000e-08 0.00000e+00
+ 2.52400e-08 0.00000e+00 2.52650e-08 6.70000e-04 2.53000e-08 0.00000e+00
+ 2.54400e-08 0.00000e+00 2.54650e-08 6.70000e-04 2.55000e-08 0.00000e+00
+ 2.56400e-08 0.00000e+00 2.56650e-08 6.70000e-04 2.57000e-08 0.00000e+00
+ 2.58400e-08 0.00000e+00 2.58650e-08 6.70000e-04 2.59000e-08 0.00000e+00
+ 2.60400e-08 0.00000e+00 2.60650e-08 6.70000e-04 2.61000e-08 0.00000e+00
+ 2.62400e-08 0.00000e+00 2.62650e-08 6.70000e-04 2.63000e-08 0.00000e+00
+ 2.64400e-08 0.00000e+00 2.64650e-08 6.70000e-04 2.65000e-08 0.00000e+00
+ 2.66400e-08 0.00000e+00 2.66650e-08 6.70000e-04 2.67000e-08 0.00000e+00
+ 2.68400e-08 0.00000e+00 2.68650e-08 6.70000e-04 2.69000e-08 0.00000e+00
+ 2.70400e-08 0.00000e+00 2.70650e-08 6.70000e-04 2.71000e-08 0.00000e+00
+ 2.72400e-08 0.00000e+00 2.72650e-08 6.70000e-04 2.73000e-08 0.00000e+00
+ 2.74400e-08 0.00000e+00 2.74650e-08 6.70000e-04 2.75000e-08 0.00000e+00
+ 2.76400e-08 0.00000e+00 2.76650e-08 6.70000e-04 2.77000e-08 0.00000e+00
+ 2.78400e-08 0.00000e+00 2.78650e-08 6.70000e-04 2.79000e-08 0.00000e+00
+ 2.80400e-08 0.00000e+00 2.80650e-08 6.70000e-04 2.81000e-08 0.00000e+00
+ 2.82400e-08 0.00000e+00 2.82650e-08 6.70000e-04 2.83000e-08 0.00000e+00
+ 2.84400e-08 0.00000e+00 2.84650e-08 6.70000e-04 2.85000e-08 0.00000e+00
+ 2.86400e-08 0.00000e+00 2.86650e-08 6.70000e-04 2.87000e-08 0.00000e+00
+ 2.88400e-08 0.00000e+00 2.88650e-08 6.70000e-04 2.89000e-08 0.00000e+00
+ 2.90400e-08 0.00000e+00 2.90650e-08 6.70000e-04 2.91000e-08 0.00000e+00
+ 2.92400e-08 0.00000e+00 2.92650e-08 6.70000e-04 2.93000e-08 0.00000e+00
+ 2.94400e-08 0.00000e+00 2.94650e-08 6.70000e-04 2.95000e-08 0.00000e+00
+ 2.96400e-08 0.00000e+00 2.96650e-08 6.70000e-04 2.97000e-08 0.00000e+00
+ 2.98400e-08 0.00000e+00 2.98650e-08 6.70000e-04 2.99000e-08 0.00000e+00
+ 3.00400e-08 0.00000e+00 3.00650e-08 6.70000e-04 3.01000e-08 0.00000e+00
+ 3.02400e-08 0.00000e+00 3.02650e-08 6.70000e-04 3.03000e-08 0.00000e+00
+ 3.04400e-08 0.00000e+00 3.04650e-08 6.70000e-04 3.05000e-08 0.00000e+00
+ 3.06400e-08 0.00000e+00 3.06650e-08 6.70000e-04 3.07000e-08 0.00000e+00
+ 3.08400e-08 0.00000e+00 3.08650e-08 6.70000e-04 3.09000e-08 0.00000e+00
+ 3.10400e-08 0.00000e+00 3.10650e-08 6.70000e-04 3.11000e-08 0.00000e+00
+ 3.12400e-08 0.00000e+00 3.12650e-08 6.70000e-04 3.13000e-08 0.00000e+00
+ 3.14400e-08 0.00000e+00 3.14650e-08 6.70000e-04 3.15000e-08 0.00000e+00
+ 3.16400e-08 0.00000e+00 3.16650e-08 6.70000e-04 3.17000e-08 0.00000e+00
+ 3.18400e-08 0.00000e+00 3.18650e-08 6.70000e-04 3.19000e-08 0.00000e+00
+ 3.20400e-08 0.00000e+00 3.20650e-08 6.70000e-04 3.21000e-08 0.00000e+00
+ 3.22400e-08 0.00000e+00 3.22650e-08 6.70000e-04 3.23000e-08 0.00000e+00
+ 3.24400e-08 0.00000e+00 3.24650e-08 6.70000e-04 3.25000e-08 0.00000e+00
+ 3.26400e-08 0.00000e+00 3.26650e-08 6.70000e-04 3.27000e-08 0.00000e+00
+ 3.28400e-08 0.00000e+00 3.28650e-08 6.70000e-04 3.29000e-08 0.00000e+00
+ 3.30400e-08 0.00000e+00 3.30650e-08 6.70000e-04 3.31000e-08 0.00000e+00
+ 3.32400e-08 0.00000e+00 3.32650e-08 6.70000e-04 3.33000e-08 0.00000e+00
+ 3.34400e-08 0.00000e+00 3.34650e-08 6.70000e-04 3.35000e-08 0.00000e+00
+ 3.36400e-08 0.00000e+00 3.36650e-08 6.70000e-04 3.37000e-08 0.00000e+00
+ 3.38400e-08 0.00000e+00 3.38650e-08 6.70000e-04 3.39000e-08 0.00000e+00
+ 3.40400e-08 0.00000e+00 3.40650e-08 6.70000e-04 3.41000e-08 0.00000e+00
+ 3.42400e-08 0.00000e+00 3.42650e-08 6.70000e-04 3.43000e-08 0.00000e+00
+ 3.44400e-08 0.00000e+00 3.44650e-08 6.70000e-04 3.45000e-08 0.00000e+00
+ 3.46400e-08 0.00000e+00 3.46650e-08 6.70000e-04 3.47000e-08 0.00000e+00
+ 3.48400e-08 0.00000e+00 3.48650e-08 6.70000e-04 3.49000e-08 0.00000e+00
+ 3.50400e-08 0.00000e+00 3.50650e-08 6.70000e-04 3.51000e-08 0.00000e+00
+ 3.52400e-08 0.00000e+00 3.52650e-08 6.70000e-04 3.53000e-08 0.00000e+00
+ 3.54400e-08 0.00000e+00 3.54650e-08 6.70000e-04 3.55000e-08 0.00000e+00
+ 3.56400e-08 0.00000e+00 3.56650e-08 6.70000e-04 3.57000e-08 0.00000e+00
+ 3.58400e-08 0.00000e+00 3.58650e-08 6.70000e-04 3.59000e-08 0.00000e+00
+ 3.60400e-08 0.00000e+00 3.60650e-08 6.70000e-04 3.61000e-08 0.00000e+00
+ 3.62400e-08 0.00000e+00 3.62650e-08 6.70000e-04 3.63000e-08 0.00000e+00
+ 3.64400e-08 0.00000e+00 3.64650e-08 6.70000e-04 3.65000e-08 0.00000e+00
+ 3.66400e-08 0.00000e+00 3.66650e-08 6.70000e-04 3.67000e-08 0.00000e+00
+ 3.68400e-08 0.00000e+00 3.68650e-08 6.70000e-04 3.69000e-08 0.00000e+00
+ 3.70400e-08 0.00000e+00 3.70650e-08 6.70000e-04 3.71000e-08 0.00000e+00
+ 3.72400e-08 0.00000e+00 3.72650e-08 6.70000e-04 3.73000e-08 0.00000e+00
+ 3.74400e-08 0.00000e+00 3.74650e-08 6.70000e-04 3.75000e-08 0.00000e+00
+ 3.76400e-08 0.00000e+00 3.76650e-08 6.70000e-04 3.77000e-08 0.00000e+00
+ 3.78400e-08 0.00000e+00 3.78650e-08 6.70000e-04 3.79000e-08 0.00000e+00
+ 3.80400e-08 0.00000e+00 3.80650e-08 6.70000e-04 3.81000e-08 0.00000e+00
+ 3.82400e-08 0.00000e+00 3.82650e-08 6.70000e-04 3.83000e-08 0.00000e+00
+ 3.84400e-08 0.00000e+00 3.84650e-08 6.70000e-04 3.85000e-08 0.00000e+00
+ 3.86400e-08 0.00000e+00 3.86650e-08 6.70000e-04 3.87000e-08 0.00000e+00
+ 3.88400e-08 0.00000e+00 3.88650e-08 6.70000e-04 3.89000e-08 0.00000e+00
+ 3.90400e-08 0.00000e+00 3.90650e-08 6.70000e-04 3.91000e-08 0.00000e+00
+ 3.92400e-08 0.00000e+00 3.92650e-08 6.70000e-04 3.93000e-08 0.00000e+00
+ 3.94400e-08 0.00000e+00 3.94650e-08 6.70000e-04 3.95000e-08 0.00000e+00
+ 3.96400e-08 0.00000e+00 3.96650e-08 6.70000e-04 3.97000e-08 0.00000e+00
+ 3.98400e-08 0.00000e+00 3.98650e-08 6.70000e-04 3.99000e-08 0.00000e+00
+ 4.00400e-08 0.00000e+00 4.00650e-08 6.70000e-04 4.01000e-08 0.00000e+00
+ 4.02400e-08 0.00000e+00 4.02650e-08 6.70000e-04 4.03000e-08 0.00000e+00
+ 4.04400e-08 0.00000e+00 4.04650e-08 6.70000e-04 4.05000e-08 0.00000e+00
+ 4.06400e-08 0.00000e+00 4.06650e-08 6.70000e-04 4.07000e-08 0.00000e+00
+ 4.08400e-08 0.00000e+00 4.08650e-08 6.70000e-04 4.09000e-08 0.00000e+00
+ 4.10400e-08 0.00000e+00 4.10650e-08 6.70000e-04 4.11000e-08 0.00000e+00
+ 4.12400e-08 0.00000e+00 4.12650e-08 6.70000e-04 4.13000e-08 0.00000e+00
+ 4.14400e-08 0.00000e+00 4.14650e-08 6.70000e-04 4.15000e-08 0.00000e+00
+ 4.16400e-08 0.00000e+00 4.16650e-08 6.70000e-04 4.17000e-08 0.00000e+00
+ 4.18400e-08 0.00000e+00 4.18650e-08 6.70000e-04 4.19000e-08 0.00000e+00
+ 4.20400e-08 0.00000e+00 4.20650e-08 6.70000e-04 4.21000e-08 0.00000e+00
+ 4.22400e-08 0.00000e+00 4.22650e-08 6.70000e-04 4.23000e-08 0.00000e+00
+ 4.24400e-08 0.00000e+00 4.24650e-08 6.70000e-04 4.25000e-08 0.00000e+00
+ 4.26400e-08 0.00000e+00 4.26650e-08 6.70000e-04 4.27000e-08 0.00000e+00
+ 4.28400e-08 0.00000e+00 4.28650e-08 6.70000e-04 4.29000e-08 0.00000e+00
+ 4.30400e-08 0.00000e+00 4.30650e-08 6.70000e-04 4.31000e-08 0.00000e+00
+ 4.32400e-08 0.00000e+00 4.32650e-08 6.70000e-04 4.33000e-08 0.00000e+00
+ 4.34400e-08 0.00000e+00 4.34650e-08 6.70000e-04 4.35000e-08 0.00000e+00
+ 4.36400e-08 0.00000e+00 4.36650e-08 6.70000e-04 4.37000e-08 0.00000e+00
+ 4.38400e-08 0.00000e+00 4.38650e-08 6.70000e-04 4.39000e-08 0.00000e+00
+ 4.40400e-08 0.00000e+00 4.40650e-08 6.70000e-04 4.41000e-08 0.00000e+00
+ 4.42400e-08 0.00000e+00 4.42650e-08 6.70000e-04 4.43000e-08 0.00000e+00
+ 4.44400e-08 0.00000e+00 4.44650e-08 6.70000e-04 4.45000e-08 0.00000e+00
+ 4.46400e-08 0.00000e+00 4.46650e-08 6.70000e-04 4.47000e-08 0.00000e+00
+ 4.48400e-08 0.00000e+00 4.48650e-08 6.70000e-04 4.49000e-08 0.00000e+00
+ 4.50400e-08 0.00000e+00 4.50650e-08 6.70000e-04 4.51000e-08 0.00000e+00
+ 4.52400e-08 0.00000e+00 4.52650e-08 6.70000e-04 4.53000e-08 0.00000e+00
+ 4.54400e-08 0.00000e+00 4.54650e-08 6.70000e-04 4.55000e-08 0.00000e+00
+ 4.56400e-08 0.00000e+00 4.56650e-08 6.70000e-04 4.57000e-08 0.00000e+00
+ 4.58400e-08 0.00000e+00 4.58650e-08 6.70000e-04 4.59000e-08 0.00000e+00
+ 4.60400e-08 0.00000e+00 4.60650e-08 6.70000e-04 4.61000e-08 0.00000e+00
+ 4.62400e-08 0.00000e+00 4.62650e-08 6.70000e-04 4.63000e-08 0.00000e+00
+ 4.64400e-08 0.00000e+00 4.64650e-08 6.70000e-04 4.65000e-08 0.00000e+00
+ 4.66400e-08 0.00000e+00 4.66650e-08 6.70000e-04 4.67000e-08 0.00000e+00
+ 4.68400e-08 0.00000e+00 4.68650e-08 6.70000e-04 4.69000e-08 0.00000e+00
+ 4.70400e-08 0.00000e+00 4.70650e-08 6.70000e-04 4.71000e-08 0.00000e+00
+ 4.72400e-08 0.00000e+00 4.72650e-08 6.70000e-04 4.73000e-08 0.00000e+00
+ 4.74400e-08 0.00000e+00 4.74650e-08 6.70000e-04 4.75000e-08 0.00000e+00
+ 4.76400e-08 0.00000e+00 4.76650e-08 6.70000e-04 4.77000e-08 0.00000e+00
+ 4.78400e-08 0.00000e+00 4.78650e-08 6.70000e-04 4.79000e-08 0.00000e+00
+ 4.80400e-08 0.00000e+00 4.80650e-08 6.70000e-04 4.81000e-08 0.00000e+00
+ 4.82400e-08 0.00000e+00 4.82650e-08 6.70000e-04 4.83000e-08 0.00000e+00
+ 4.84400e-08 0.00000e+00 4.84650e-08 6.70000e-04 4.85000e-08 0.00000e+00
+ 4.86400e-08 0.00000e+00 4.86650e-08 6.70000e-04 4.87000e-08 0.00000e+00
+ 4.88400e-08 0.00000e+00 4.88650e-08 6.70000e-04 4.89000e-08 0.00000e+00
+ 4.90400e-08 0.00000e+00 4.90650e-08 6.70000e-04 4.91000e-08 0.00000e+00
+ 4.92400e-08 0.00000e+00 4.92650e-08 6.70000e-04 4.93000e-08 0.00000e+00
+ 4.94400e-08 0.00000e+00 4.94650e-08 6.70000e-04 4.95000e-08 0.00000e+00
+ 4.96400e-08 0.00000e+00 4.96650e-08 6.70000e-04 4.97000e-08 0.00000e+00
+ 4.98400e-08 0.00000e+00 4.98650e-08 6.70000e-04 4.99000e-08 0.00000e+00
+ 5.00400e-08 0.00000e+00 5.00650e-08 6.70000e-04 5.01000e-08 0.00000e+00
+ 5.02400e-08 0.00000e+00 5.02650e-08 6.70000e-04 5.03000e-08 0.00000e+00
+ 5.04400e-08 0.00000e+00 5.04650e-08 6.70000e-04 5.05000e-08 0.00000e+00
+ 5.06400e-08 0.00000e+00 5.06650e-08 6.70000e-04 5.07000e-08 0.00000e+00
+ 5.08400e-08 0.00000e+00 5.08650e-08 6.70000e-04 5.09000e-08 0.00000e+00
+ 5.10400e-08 0.00000e+00 5.10650e-08 6.70000e-04 5.11000e-08 0.00000e+00
+ 5.12400e-08 0.00000e+00 5.12650e-08 6.70000e-04 5.13000e-08 0.00000e+00
+ 5.14400e-08 0.00000e+00 5.14650e-08 6.70000e-04 5.15000e-08 0.00000e+00
+ 5.16400e-08 0.00000e+00 5.16650e-08 6.70000e-04 5.17000e-08 0.00000e+00
+ 5.18400e-08 0.00000e+00 5.18650e-08 6.70000e-04 5.19000e-08 0.00000e+00
+ 5.20400e-08 0.00000e+00 5.20650e-08 6.70000e-04 5.21000e-08 0.00000e+00
+ 5.22400e-08 0.00000e+00 5.22650e-08 6.70000e-04 5.23000e-08 0.00000e+00
+ 5.24400e-08 0.00000e+00 5.24650e-08 6.70000e-04 5.25000e-08 0.00000e+00
+ 5.26400e-08 0.00000e+00 5.26650e-08 6.70000e-04 5.27000e-08 0.00000e+00
+ 5.28400e-08 0.00000e+00 5.28650e-08 6.70000e-04 5.29000e-08 0.00000e+00
+ 5.30400e-08 0.00000e+00 5.30650e-08 6.70000e-04 5.31000e-08 0.00000e+00
+ 5.32400e-08 0.00000e+00 5.32650e-08 6.70000e-04 5.33000e-08 0.00000e+00
+ 5.34400e-08 0.00000e+00 5.34650e-08 6.70000e-04 5.35000e-08 0.00000e+00
+ 5.36400e-08 0.00000e+00 5.36650e-08 6.70000e-04 5.37000e-08 0.00000e+00
+ 5.38400e-08 0.00000e+00 5.38650e-08 6.70000e-04 5.39000e-08 0.00000e+00
+ 5.40400e-08 0.00000e+00 5.40650e-08 6.70000e-04 5.41000e-08 0.00000e+00
+ 5.42400e-08 0.00000e+00 5.42650e-08 6.70000e-04 5.43000e-08 0.00000e+00
+ 5.44400e-08 0.00000e+00 5.44650e-08 6.70000e-04 5.45000e-08 0.00000e+00
+ 5.46400e-08 0.00000e+00 5.46650e-08 6.70000e-04 5.47000e-08 0.00000e+00
+ 5.48400e-08 0.00000e+00 5.48650e-08 6.70000e-04 5.49000e-08 0.00000e+00
+ 5.50400e-08 0.00000e+00 5.50650e-08 6.70000e-04 5.51000e-08 0.00000e+00
+ 5.52400e-08 0.00000e+00 5.52650e-08 6.70000e-04 5.53000e-08 0.00000e+00
+ 5.54400e-08 0.00000e+00 5.54650e-08 6.70000e-04 5.55000e-08 0.00000e+00
+ 5.56400e-08 0.00000e+00 5.56650e-08 6.70000e-04 5.57000e-08 0.00000e+00
+ 5.58400e-08 0.00000e+00 5.58650e-08 6.70000e-04 5.59000e-08 0.00000e+00
+ 5.60400e-08 0.00000e+00 5.60650e-08 6.70000e-04 5.61000e-08 0.00000e+00
+ 5.62400e-08 0.00000e+00 5.62650e-08 6.70000e-04 5.63000e-08 0.00000e+00
+ 5.64400e-08 0.00000e+00 5.64650e-08 6.70000e-04 5.65000e-08 0.00000e+00
+ 5.66400e-08 0.00000e+00 5.66650e-08 6.70000e-04 5.67000e-08 0.00000e+00
+ 5.68400e-08 0.00000e+00 5.68650e-08 6.70000e-04 5.69000e-08 0.00000e+00
+ 5.70400e-08 0.00000e+00 5.70650e-08 6.70000e-04 5.71000e-08 0.00000e+00
+ 5.72400e-08 0.00000e+00 5.72650e-08 6.70000e-04 5.73000e-08 0.00000e+00
+ 5.74400e-08 0.00000e+00 5.74650e-08 6.70000e-04 5.75000e-08 0.00000e+00
+ 5.76400e-08 0.00000e+00 5.76650e-08 6.70000e-04 5.77000e-08 0.00000e+00
+ 5.78400e-08 0.00000e+00 5.78650e-08 6.70000e-04 5.79000e-08 0.00000e+00
+ 5.80400e-08 0.00000e+00 5.80650e-08 6.70000e-04 5.81000e-08 0.00000e+00
+ 5.82400e-08 0.00000e+00 5.82650e-08 6.70000e-04 5.83000e-08 0.00000e+00
+ 5.84400e-08 0.00000e+00 5.84650e-08 6.70000e-04 5.85000e-08 0.00000e+00
+ 5.86400e-08 0.00000e+00 5.86650e-08 6.70000e-04 5.87000e-08 0.00000e+00
+ 5.88400e-08 0.00000e+00 5.88650e-08 6.70000e-04 5.89000e-08 0.00000e+00
+ 5.90400e-08 0.00000e+00 5.90650e-08 6.70000e-04 5.91000e-08 0.00000e+00
+ 5.92400e-08 0.00000e+00 5.92650e-08 6.70000e-04 5.93000e-08 0.00000e+00
+ 5.94400e-08 0.00000e+00 5.94650e-08 6.70000e-04 5.95000e-08 0.00000e+00
+ 5.96400e-08 0.00000e+00 5.96650e-08 6.70000e-04 5.97000e-08 0.00000e+00
+ 5.98400e-08 0.00000e+00 5.98650e-08 6.70000e-04 5.99000e-08 0.00000e+00
+ 6.00400e-08 0.00000e+00 6.00650e-08 6.70000e-04 6.01000e-08 0.00000e+00
+ 6.02400e-08 0.00000e+00 6.02650e-08 6.70000e-04 6.03000e-08 0.00000e+00
+ 6.04400e-08 0.00000e+00 6.04650e-08 6.70000e-04 6.05000e-08 0.00000e+00
+ 6.06400e-08 0.00000e+00 6.06650e-08 6.70000e-04 6.07000e-08 0.00000e+00
+ 6.08400e-08 0.00000e+00 6.08650e-08 6.70000e-04 6.09000e-08 0.00000e+00
+ 6.10400e-08 0.00000e+00 6.10650e-08 6.70000e-04 6.11000e-08 0.00000e+00
+ 6.12400e-08 0.00000e+00 6.12650e-08 6.70000e-04 6.13000e-08 0.00000e+00
+ 6.14400e-08 0.00000e+00 6.14650e-08 6.70000e-04 6.15000e-08 0.00000e+00
+ 6.16400e-08 0.00000e+00 6.16650e-08 6.70000e-04 6.17000e-08 0.00000e+00
+ 6.18400e-08 0.00000e+00 6.18650e-08 6.70000e-04 6.19000e-08 0.00000e+00
+ 6.20400e-08 0.00000e+00 6.20650e-08 6.70000e-04 6.21000e-08 0.00000e+00
+ 6.22400e-08 0.00000e+00 6.22650e-08 6.70000e-04 6.23000e-08 0.00000e+00
+ 6.24400e-08 0.00000e+00 6.24650e-08 6.70000e-04 6.25000e-08 0.00000e+00
+ 6.26400e-08 0.00000e+00 6.26650e-08 6.70000e-04 6.27000e-08 0.00000e+00
+ 6.28400e-08 0.00000e+00 6.28650e-08 6.70000e-04 6.29000e-08 0.00000e+00
+ 6.30400e-08 0.00000e+00 6.30650e-08 6.70000e-04 6.31000e-08 0.00000e+00
+ 6.32400e-08 0.00000e+00 6.32650e-08 6.70000e-04 6.33000e-08 0.00000e+00
+ 6.34400e-08 0.00000e+00 6.34650e-08 6.70000e-04 6.35000e-08 0.00000e+00
+ 6.36400e-08 0.00000e+00 6.36650e-08 6.70000e-04 6.37000e-08 0.00000e+00
+ 6.38400e-08 0.00000e+00 6.38650e-08 6.70000e-04 6.39000e-08 0.00000e+00
+ 6.40400e-08 0.00000e+00 6.40650e-08 6.70000e-04 6.41000e-08 0.00000e+00
+ 6.42400e-08 0.00000e+00 6.42650e-08 6.70000e-04 6.43000e-08 0.00000e+00
+ 6.44400e-08 0.00000e+00 6.44650e-08 6.70000e-04 6.45000e-08 0.00000e+00
+ 6.46400e-08 0.00000e+00 6.46650e-08 6.70000e-04 6.47000e-08 0.00000e+00
+ 6.48400e-08 0.00000e+00 6.48650e-08 6.70000e-04 6.49000e-08 0.00000e+00
+ 6.50400e-08 0.00000e+00 6.50650e-08 6.70000e-04 6.51000e-08 0.00000e+00
+ 6.52400e-08 0.00000e+00 6.52650e-08 6.70000e-04 6.53000e-08 0.00000e+00
+ 6.54400e-08 0.00000e+00 6.54650e-08 6.70000e-04 6.55000e-08 0.00000e+00
+ 6.56400e-08 0.00000e+00 6.56650e-08 6.70000e-04 6.57000e-08 0.00000e+00
+ 6.58400e-08 0.00000e+00 6.58650e-08 6.70000e-04 6.59000e-08 0.00000e+00
+ 6.60400e-08 0.00000e+00 6.60650e-08 6.70000e-04 6.61000e-08 0.00000e+00
+ 6.62400e-08 0.00000e+00 6.62650e-08 6.70000e-04 6.63000e-08 0.00000e+00
+ 6.64400e-08 0.00000e+00 6.64650e-08 6.70000e-04 6.65000e-08 0.00000e+00
+ 6.66400e-08 0.00000e+00 6.66650e-08 6.70000e-04 6.67000e-08 0.00000e+00
+ 6.68400e-08 0.00000e+00 6.68650e-08 6.70000e-04 6.69000e-08 0.00000e+00
+ 6.70400e-08 0.00000e+00 6.70650e-08 6.70000e-04 6.71000e-08 0.00000e+00
+ 6.72400e-08 0.00000e+00 6.72650e-08 6.70000e-04 6.73000e-08 0.00000e+00
+ 6.74400e-08 0.00000e+00 6.74650e-08 6.70000e-04 6.75000e-08 0.00000e+00
+ 6.76400e-08 0.00000e+00 6.76650e-08 6.70000e-04 6.77000e-08 0.00000e+00
+ 6.78400e-08 0.00000e+00 6.78650e-08 6.70000e-04 6.79000e-08 0.00000e+00
+ 6.80400e-08 0.00000e+00 6.80650e-08 6.70000e-04 6.81000e-08 0.00000e+00
+ 6.82400e-08 0.00000e+00 6.82650e-08 6.70000e-04 6.83000e-08 0.00000e+00
+ 6.84400e-08 0.00000e+00 6.84650e-08 6.70000e-04 6.85000e-08 0.00000e+00
+ 6.86400e-08 0.00000e+00 6.86650e-08 6.70000e-04 6.87000e-08 0.00000e+00
+ 6.88400e-08 0.00000e+00 6.88650e-08 6.70000e-04 6.89000e-08 0.00000e+00
+ 6.90400e-08 0.00000e+00 6.90650e-08 6.70000e-04 6.91000e-08 0.00000e+00
+ 6.92400e-08 0.00000e+00 6.92650e-08 6.70000e-04 6.93000e-08 0.00000e+00
+ 6.94400e-08 0.00000e+00 6.94650e-08 6.70000e-04 6.95000e-08 0.00000e+00
+ 6.96400e-08 0.00000e+00 6.96650e-08 6.70000e-04 6.97000e-08 0.00000e+00
+ 6.98400e-08 0.00000e+00 6.98650e-08 6.70000e-04 6.99000e-08 0.00000e+00
+ 7.00400e-08 0.00000e+00 7.00650e-08 6.70000e-04 7.01000e-08 0.00000e+00
+ 7.02400e-08 0.00000e+00 7.02650e-08 6.70000e-04 7.03000e-08 0.00000e+00
+ 7.04400e-08 0.00000e+00 7.04650e-08 6.70000e-04 7.05000e-08 0.00000e+00
+ 7.06400e-08 0.00000e+00 7.06650e-08 6.70000e-04 7.07000e-08 0.00000e+00
+ 7.08400e-08 0.00000e+00 7.08650e-08 6.70000e-04 7.09000e-08 0.00000e+00
+ 7.10400e-08 0.00000e+00 7.10650e-08 6.70000e-04 7.11000e-08 0.00000e+00
+ 7.12400e-08 0.00000e+00 7.12650e-08 6.70000e-04 7.13000e-08 0.00000e+00
+ 7.14400e-08 0.00000e+00 7.14650e-08 6.70000e-04 7.15000e-08 0.00000e+00
+ 7.16400e-08 0.00000e+00 7.16650e-08 6.70000e-04 7.17000e-08 0.00000e+00
+ 7.18400e-08 0.00000e+00 7.18650e-08 6.70000e-04 7.19000e-08 0.00000e+00
+ 7.20400e-08 0.00000e+00 7.20650e-08 6.70000e-04 7.21000e-08 0.00000e+00
+ 7.22400e-08 0.00000e+00 7.22650e-08 6.70000e-04 7.23000e-08 0.00000e+00
+ 7.24400e-08 0.00000e+00 7.24650e-08 6.70000e-04 7.25000e-08 0.00000e+00
+ 7.26400e-08 0.00000e+00 7.26650e-08 6.70000e-04 7.27000e-08 0.00000e+00
+ 7.28400e-08 0.00000e+00 7.28650e-08 6.70000e-04 7.29000e-08 0.00000e+00
+ 7.30400e-08 0.00000e+00 7.30650e-08 6.70000e-04 7.31000e-08 0.00000e+00
+ 7.32400e-08 0.00000e+00 7.32650e-08 6.70000e-04 7.33000e-08 0.00000e+00
+ 7.34400e-08 0.00000e+00 7.34650e-08 6.70000e-04 7.35000e-08 0.00000e+00
+ 7.36400e-08 0.00000e+00 7.36650e-08 6.70000e-04 7.37000e-08 0.00000e+00
+ 7.38400e-08 0.00000e+00 7.38650e-08 6.70000e-04 7.39000e-08 0.00000e+00
+ 7.40400e-08 0.00000e+00 7.40650e-08 6.70000e-04 7.41000e-08 0.00000e+00
+ 7.42400e-08 0.00000e+00 7.42650e-08 6.70000e-04 7.43000e-08 0.00000e+00
+ 7.44400e-08 0.00000e+00 7.44650e-08 6.70000e-04 7.45000e-08 0.00000e+00
+ 7.46400e-08 0.00000e+00 7.46650e-08 6.70000e-04 7.47000e-08 0.00000e+00
+ 7.48400e-08 0.00000e+00 7.48650e-08 6.70000e-04 7.49000e-08 0.00000e+00
+ 7.50400e-08 0.00000e+00 7.50650e-08 6.70000e-04 7.51000e-08 0.00000e+00
+ 7.52400e-08 0.00000e+00 7.52650e-08 6.70000e-04 7.53000e-08 0.00000e+00
+ 7.54400e-08 0.00000e+00 7.54650e-08 6.70000e-04 7.55000e-08 0.00000e+00
+ 7.56400e-08 0.00000e+00 7.56650e-08 6.70000e-04 7.57000e-08 0.00000e+00
+ 7.58400e-08 0.00000e+00 7.58650e-08 6.70000e-04 7.59000e-08 0.00000e+00
+ 7.60400e-08 0.00000e+00 7.60650e-08 6.70000e-04 7.61000e-08 0.00000e+00
+ 7.62400e-08 0.00000e+00 7.62650e-08 6.70000e-04 7.63000e-08 0.00000e+00
+ 7.64400e-08 0.00000e+00 7.64650e-08 6.70000e-04 7.65000e-08 0.00000e+00
+ 7.66400e-08 0.00000e+00 7.66650e-08 6.70000e-04 7.67000e-08 0.00000e+00
+ 7.68400e-08 0.00000e+00 7.68650e-08 6.70000e-04 7.69000e-08 0.00000e+00
+ 7.70400e-08 0.00000e+00 7.70650e-08 6.70000e-04 7.71000e-08 0.00000e+00
+ 7.72400e-08 0.00000e+00 7.72650e-08 6.70000e-04 7.73000e-08 0.00000e+00
+ 7.74400e-08 0.00000e+00 7.74650e-08 6.70000e-04 7.75000e-08 0.00000e+00
+ 7.76400e-08 0.00000e+00 7.76650e-08 6.70000e-04 7.77000e-08 0.00000e+00
+ 7.78400e-08 0.00000e+00 7.78650e-08 6.70000e-04 7.79000e-08 0.00000e+00
+ 7.80400e-08 0.00000e+00 7.80650e-08 6.70000e-04 7.81000e-08 0.00000e+00
+ 7.82400e-08 0.00000e+00 7.82650e-08 6.70000e-04 7.83000e-08 0.00000e+00
+ 7.84400e-08 0.00000e+00 7.84650e-08 6.70000e-04 7.85000e-08 0.00000e+00
+ 7.86400e-08 0.00000e+00 7.86650e-08 6.70000e-04 7.87000e-08 0.00000e+00
+ 7.88400e-08 0.00000e+00 7.88650e-08 6.70000e-04 7.89000e-08 0.00000e+00
+ 7.90400e-08 0.00000e+00 7.90650e-08 6.70000e-04 7.91000e-08 0.00000e+00
+ 7.92400e-08 0.00000e+00 7.92650e-08 6.70000e-04 7.93000e-08 0.00000e+00
+ 7.94400e-08 0.00000e+00 7.94650e-08 6.70000e-04 7.95000e-08 0.00000e+00
+ 7.96400e-08 0.00000e+00 7.96650e-08 6.70000e-04 7.97000e-08 0.00000e+00
+ 7.98400e-08 0.00000e+00 7.98650e-08 6.70000e-04 7.99000e-08 0.00000e+00
+ 8.00400e-08 0.00000e+00 8.00650e-08 6.70000e-04 8.01000e-08 0.00000e+00
+ 8.02400e-08 0.00000e+00 8.02650e-08 6.70000e-04 8.03000e-08 0.00000e+00
+ 8.04400e-08 0.00000e+00 8.04650e-08 6.70000e-04 8.05000e-08 0.00000e+00
+ 8.06400e-08 0.00000e+00 8.06650e-08 6.70000e-04 8.07000e-08 0.00000e+00
+ 8.08400e-08 0.00000e+00 8.08650e-08 6.70000e-04 8.09000e-08 0.00000e+00
+ 8.10400e-08 0.00000e+00 8.10650e-08 6.70000e-04 8.11000e-08 0.00000e+00
+ 8.12400e-08 0.00000e+00 8.12650e-08 6.70000e-04 8.13000e-08 0.00000e+00
+ 8.14400e-08 0.00000e+00 8.14650e-08 6.70000e-04 8.15000e-08 0.00000e+00
+ 8.16400e-08 0.00000e+00 8.16650e-08 6.70000e-04 8.17000e-08 0.00000e+00
+ 8.18400e-08 0.00000e+00 8.18650e-08 6.70000e-04 8.19000e-08 0.00000e+00
+ 8.20400e-08 0.00000e+00 8.20650e-08 6.70000e-04 8.21000e-08 0.00000e+00
+ 8.22400e-08 0.00000e+00 8.22650e-08 6.70000e-04 8.23000e-08 0.00000e+00
+ 8.24400e-08 0.00000e+00 8.24650e-08 6.70000e-04 8.25000e-08 0.00000e+00
+ 8.26400e-08 0.00000e+00 8.26650e-08 6.70000e-04 8.27000e-08 0.00000e+00
+ 8.28400e-08 0.00000e+00 8.28650e-08 6.70000e-04 8.29000e-08 0.00000e+00
+ 8.30400e-08 0.00000e+00 8.30650e-08 6.70000e-04 8.31000e-08 0.00000e+00
+ 8.32400e-08 0.00000e+00 8.32650e-08 6.70000e-04 8.33000e-08 0.00000e+00
+ 8.34400e-08 0.00000e+00 8.34650e-08 6.70000e-04 8.35000e-08 0.00000e+00
+ 8.36400e-08 0.00000e+00 8.36650e-08 6.70000e-04 8.37000e-08 0.00000e+00
+ 8.38400e-08 0.00000e+00 8.38650e-08 6.70000e-04 8.39000e-08 0.00000e+00
+ 8.40400e-08 0.00000e+00 8.40650e-08 6.70000e-04 8.41000e-08 0.00000e+00
+ 8.42400e-08 0.00000e+00 8.42650e-08 6.70000e-04 8.43000e-08 0.00000e+00
+ 8.44400e-08 0.00000e+00 8.44650e-08 6.70000e-04 8.45000e-08 0.00000e+00
+ 8.46400e-08 0.00000e+00 8.46650e-08 6.70000e-04 8.47000e-08 0.00000e+00
+ 8.48400e-08 0.00000e+00 8.48650e-08 6.70000e-04 8.49000e-08 0.00000e+00
+ 8.50400e-08 0.00000e+00 8.50650e-08 6.70000e-04 8.51000e-08 0.00000e+00
+ 8.52400e-08 0.00000e+00 8.52650e-08 6.70000e-04 8.53000e-08 0.00000e+00
+ 8.54400e-08 0.00000e+00 8.54650e-08 6.70000e-04 8.55000e-08 0.00000e+00
+ 8.56400e-08 0.00000e+00 8.56650e-08 6.70000e-04 8.57000e-08 0.00000e+00
+ 8.58400e-08 0.00000e+00 8.58650e-08 6.70000e-04 8.59000e-08 0.00000e+00
+ 8.60400e-08 0.00000e+00 8.60650e-08 6.70000e-04 8.61000e-08 0.00000e+00
+ 8.62400e-08 0.00000e+00 8.62650e-08 6.70000e-04 8.63000e-08 0.00000e+00
+ 8.64400e-08 0.00000e+00 8.64650e-08 6.70000e-04 8.65000e-08 0.00000e+00
+ 8.66400e-08 0.00000e+00 8.66650e-08 6.70000e-04 8.67000e-08 0.00000e+00
+ 8.68400e-08 0.00000e+00 8.68650e-08 6.70000e-04 8.69000e-08 0.00000e+00
+ 8.70400e-08 0.00000e+00 8.70650e-08 6.70000e-04 8.71000e-08 0.00000e+00
+ 8.72400e-08 0.00000e+00 8.72650e-08 6.70000e-04 8.73000e-08 0.00000e+00
+ 8.74400e-08 0.00000e+00 8.74650e-08 6.70000e-04 8.75000e-08 0.00000e+00
+ 8.76400e-08 0.00000e+00 8.76650e-08 6.70000e-04 8.77000e-08 0.00000e+00
+ 8.78400e-08 0.00000e+00 8.78650e-08 6.70000e-04 8.79000e-08 0.00000e+00
+ 8.80400e-08 0.00000e+00 8.80650e-08 6.70000e-04 8.81000e-08 0.00000e+00
+ 8.82400e-08 0.00000e+00 8.82650e-08 6.70000e-04 8.83000e-08 0.00000e+00
+ 8.84400e-08 0.00000e+00 8.84650e-08 6.70000e-04 8.85000e-08 0.00000e+00
+ 8.86400e-08 0.00000e+00 8.86650e-08 6.70000e-04 8.87000e-08 0.00000e+00
+ 8.88400e-08 0.00000e+00 8.88650e-08 6.70000e-04 8.89000e-08 0.00000e+00
+ 8.90400e-08 0.00000e+00 8.90650e-08 6.70000e-04 8.91000e-08 0.00000e+00
+ 8.92400e-08 0.00000e+00 8.92650e-08 6.70000e-04 8.93000e-08 0.00000e+00
+ 8.94400e-08 0.00000e+00 8.94650e-08 6.70000e-04 8.95000e-08 0.00000e+00
+ 8.96400e-08 0.00000e+00 8.96650e-08 6.70000e-04 8.97000e-08 0.00000e+00
+ 8.98400e-08 0.00000e+00 8.98650e-08 6.70000e-04 8.99000e-08 0.00000e+00
+ 9.00400e-08 0.00000e+00 9.00650e-08 6.70000e-04 9.01000e-08 0.00000e+00
+ 9.02400e-08 0.00000e+00 9.02650e-08 6.70000e-04 9.03000e-08 0.00000e+00
+ 9.04400e-08 0.00000e+00 9.04650e-08 6.70000e-04 9.05000e-08 0.00000e+00
+ 9.06400e-08 0.00000e+00 9.06650e-08 6.70000e-04 9.07000e-08 0.00000e+00
+ 9.08400e-08 0.00000e+00 9.08650e-08 6.70000e-04 9.09000e-08 0.00000e+00
+ 9.10400e-08 0.00000e+00 9.10650e-08 6.70000e-04 9.11000e-08 0.00000e+00
+ 9.12400e-08 0.00000e+00 9.12650e-08 6.70000e-04 9.13000e-08 0.00000e+00
+ 9.14400e-08 0.00000e+00 9.14650e-08 6.70000e-04 9.15000e-08 0.00000e+00
+ 9.16400e-08 0.00000e+00 9.16650e-08 6.70000e-04 9.17000e-08 0.00000e+00
+ 9.18400e-08 0.00000e+00 9.18650e-08 6.70000e-04 9.19000e-08 0.00000e+00
+ 9.20400e-08 0.00000e+00 9.20650e-08 6.70000e-04 9.21000e-08 0.00000e+00
+ 9.22400e-08 0.00000e+00 9.22650e-08 6.70000e-04 9.23000e-08 0.00000e+00
+ 9.24400e-08 0.00000e+00 9.24650e-08 6.70000e-04 9.25000e-08 0.00000e+00
+ 9.26400e-08 0.00000e+00 9.26650e-08 6.70000e-04 9.27000e-08 0.00000e+00
+ 9.28400e-08 0.00000e+00 9.28650e-08 6.70000e-04 9.29000e-08 0.00000e+00
+ 9.30400e-08 0.00000e+00 9.30650e-08 6.70000e-04 9.31000e-08 0.00000e+00
+ 9.32400e-08 0.00000e+00 9.32650e-08 6.70000e-04 9.33000e-08 0.00000e+00
+ 9.34400e-08 0.00000e+00 9.34650e-08 6.70000e-04 9.35000e-08 0.00000e+00
+ 9.36400e-08 0.00000e+00 9.36650e-08 6.70000e-04 9.37000e-08 0.00000e+00
+ 9.38400e-08 0.00000e+00 9.38650e-08 6.70000e-04 9.39000e-08 0.00000e+00
+ 9.40400e-08 0.00000e+00 9.40650e-08 6.70000e-04 9.41000e-08 0.00000e+00
+ 9.42400e-08 0.00000e+00 9.42650e-08 6.70000e-04 9.43000e-08 0.00000e+00
+ 9.44400e-08 0.00000e+00 9.44650e-08 6.70000e-04 9.45000e-08 0.00000e+00
+ 9.46400e-08 0.00000e+00 9.46650e-08 6.70000e-04 9.47000e-08 0.00000e+00
+ 9.48400e-08 0.00000e+00 9.48650e-08 6.70000e-04 9.49000e-08 0.00000e+00
+ 9.50400e-08 0.00000e+00 9.50650e-08 6.70000e-04 9.51000e-08 0.00000e+00
+ 9.52400e-08 0.00000e+00 9.52650e-08 6.70000e-04 9.53000e-08 0.00000e+00
+ 9.54400e-08 0.00000e+00 9.54650e-08 6.70000e-04 9.55000e-08 0.00000e+00
+ 9.56400e-08 0.00000e+00 9.56650e-08 6.70000e-04 9.57000e-08 0.00000e+00
+ 9.58400e-08 0.00000e+00 9.58650e-08 6.70000e-04 9.59000e-08 0.00000e+00
+ 9.60400e-08 0.00000e+00 9.60650e-08 6.70000e-04 9.61000e-08 0.00000e+00
+ 9.62400e-08 0.00000e+00 9.62650e-08 6.70000e-04 9.63000e-08 0.00000e+00
+ 9.64400e-08 0.00000e+00 9.64650e-08 6.70000e-04 9.65000e-08 0.00000e+00
+ 9.66400e-08 0.00000e+00 9.66650e-08 6.70000e-04 9.67000e-08 0.00000e+00
+ 9.68400e-08 0.00000e+00 9.68650e-08 6.70000e-04 9.69000e-08 0.00000e+00
+ 9.70400e-08 0.00000e+00 9.70650e-08 6.70000e-04 9.71000e-08 0.00000e+00
+ 9.72400e-08 0.00000e+00 9.72650e-08 6.70000e-04 9.73000e-08 0.00000e+00
+ 9.74400e-08 0.00000e+00 9.74650e-08 6.70000e-04 9.75000e-08 0.00000e+00
+ 9.76400e-08 0.00000e+00 9.76650e-08 6.70000e-04 9.77000e-08 0.00000e+00
+ 9.78400e-08 0.00000e+00 9.78650e-08 6.70000e-04 9.79000e-08 0.00000e+00
+ 9.80400e-08 0.00000e+00 9.80650e-08 6.70000e-04 9.81000e-08 0.00000e+00
+ 9.82400e-08 0.00000e+00 9.82650e-08 6.70000e-04 9.83000e-08 0.00000e+00
+ 9.84400e-08 0.00000e+00 9.84650e-08 6.70000e-04 9.85000e-08 0.00000e+00
+ 9.86400e-08 0.00000e+00 9.86650e-08 6.70000e-04 9.87000e-08 0.00000e+00
+ 9.88400e-08 0.00000e+00 9.88650e-08 6.70000e-04 9.89000e-08 0.00000e+00
+ 9.90400e-08 0.00000e+00 9.90650e-08 6.70000e-04 9.91000e-08 0.00000e+00
+ 9.92400e-08 0.00000e+00 9.92650e-08 6.70000e-04 9.93000e-08 0.00000e+00
+ 9.94400e-08 0.00000e+00 9.94650e-08 6.70000e-04 9.95000e-08 0.00000e+00
+ 9.96400e-08 0.00000e+00 9.96650e-08 6.70000e-04 9.97000e-08 0.00000e+00
+ 9.98400e-08 0.00000e+00 9.98650e-08 6.70000e-04 9.99000e-08 0.00000e+00
+ 1.00040e-07 0.00000e+00 1.00065e-07 6.70000e-04 1.00100e-07 0.00000e+00
+ 1.00240e-07 0.00000e+00 1.00265e-07 6.70000e-04 1.00300e-07 0.00000e+00
+ 1.00440e-07 0.00000e+00 1.00465e-07 6.70000e-04 1.00500e-07 0.00000e+00)

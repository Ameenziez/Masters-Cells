#SPLIT INTO 8 SFQ PULSES
.subckt MULTISPLIT IN SPLIT7 SPLIT8 SPLIT9 SPLIT10 SPLIT11 SPLIT12 SPLIT13 SPLIT14

#INITIAL SPLITS
XSPLIT0 LSmitll_SPLITT IN split1 split2
XSPLIT1 LSmitll_SPLITT SPLIT1 split3 split4
XSPLIT2 LSmitll_SPLITT SPLIT2 split5 split6
#use these AS OUTPUT SFQS
XSPLIT3 LSmitll_SPLITT SPLIT3 split7 split8
XSPLIT4 LSmitll_SPLITT SPLIT4 split9 split10
XSPLIT5 LSmitll_SPLITT SPLIT5 split11 split12
XSPLIT6 LSmitll_SPLITT SPLIT6 split13 split14

.ENDS MULTISPLIT
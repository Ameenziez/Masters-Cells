#works well!
#got the data to propagate
.include LSmitll_DCSFQ_PTLTX_v1p5.cir
.include LSmitll_bufft_v1p5.cir
.include LSmitll_PTLRX_SFQDC_v1p5.cir
.include LSmitll_SPLITT_v1p5.cir
.INCLUDE LSMITLL_JTLT_V1P5.CIR
.INCLUDE LSMITLL_MERGET_V1P5.CIR
.include storeedit.cir
.INCLUDE COMPONENTSEDIT.CIR
.INCLUDE COMP3.CIR
.INCLUDE COMP4.CIR
.INCLUDE COMP5.CIR
.INCLUDE COMP6.CIR
.include conv.cir
.INCLUDE synapsenext2.CIR
.INCLUDE DCPULSER.CIR
.INCLUDE MULTISPLIT.CIR
.include transmit.cir
.INCLUDE DELAY7.CIR
.INCLUDE AND.CIR
.INCLUDE AND3.CIR
.INCLUDE OR3.CIR
.include PERCEPTRON.CIR
.include PERCEPTRON2.CIR
.include CONVINTERFACE.cir


# TRY SHIFTING CLK OF OUTPUT BACK A BIT...

.tran 1ps 25000PS 0ps 1p
#MLP:
#D=Oi.T + Oi.!Oj + T.!Oj 

#setup circuitry
VAC1   A1   0   SIN(0 723mV 10GHz 200Ps 0)
RAC1   A1   A2   1000
LAC1   A2   A3   0.1p
VAC2   B1   0   SIN(0 723mV 10GHz 175.0ps 0)
RAC2   B1   B2   1000
LAC2   B2   B3   0.1p
VDC    DC1   0   pwl(0 0 20p 1023mV)
RDC    DC1   DC2   1000
LDC    DC2   DC3  0.1p
VDCconv    DCc1   0   PWL(0ps 0mV 20ps 1023mV 1.881e-08 1023mV )
RDCconv    DCc1   DCc2  640
LDCconv    DCc2   DCc3   0.1p




#SECOND LAYER SYNAPSE 1
#IINITAL21 0 INITIAL21 PWL( 0 0 20P flx21*2*-22.6U 5000p flx21*2*-22.6U 5001p 0)
IINITAL21 0 INITIAL21 PWL( 0 0 20P flx21*2*-22.6U 5000p flx21*2*-22.6U)

XSTORE21 BISTORE SFQOUTPLUS21 SFQOUTMINUS21 WEIGHTL21 WEIGHTR21


#NEXT LAYER BIAS
#Iactualsynbias21 0 ACTUALSYNB21x PWL(0 0 640P 0 665P 670U 700P 0 840P 0 865P 670U 900P 0  1040P 0 1065P 670U 1100P 0 1240P 0 1265P 670U 1300P 0  )
LSYNB21 ACTUALSYNB21x ACTUALSYNB21 1p  
KSYNB21 LSYNB21 LSYNADJUSTB21 0.3
#KSYNB21 LSYNB21 LSYNADJUSTB21 -0.3
LSYNADJUSTB21 0 ADJUSTB21 5P 

#SPLIT TARGET BETWEEN 2 NEURONS
LTARGET1 TARGET0 TARGET1 1p
LTARGET2 TARGET0 TARGET2 1p

#SPLIT INPUTS BETWEEN 2 NEURONS
LINPUT1 IN1 INPUT11 1P
LINPUT2 IN1 INPUT12 1P
LINPUT3 IN2 INPUT13 1P
LINPUT4 IN2 INPUT14 1P
LINPUTBIAS11 INB11 INPUTB12 1P
LINPUTBIAS12 INB11 INPUTB13 1P


#IINITALB21 0 INITIALB21 PWL( 0 0 20P flxb21*2*22.6U 5000p flxb21*2*22.6U 5001p 0)
IINITALB21 0 INITIALB21 PWL( 0 0 20P flxb21*2*22.6U 5000p flxb21*2*22.6U)

XSTOREB21 BISTORE SFQOUTPLUSB21 SFQOUTMINUSB21 WEIGHTLB21 WEIGHTRB21

X21 SYNAPSEfastestnext2 OUTPUTAXON DOUT22 DOUT21  WEIGHTL21 WEIGHTR21 INITIAL21
XB21 SYNAPSEfastestnext2 ACTUALSYNB21  0 DOUT23   WEIGHTLB21 WEIGHTRB21 INITIALB21

.param flx11 = -2
.param flx12 = 2
.param flx13 = 3
.param flx14 = 0
.param flxb11 = 1
.param flxb12 = -1
.param flx21 = -4
.param flx22 = 3
.param flxb21 = 0


IINITAL11 0 INITIAL11 PWL( 0 0 20P -22U*2*flx11 5000p -22U*2*flx11 5001p 0)
IINITAL12 0 INITIAL12 PWL( 0 0 20P -22u*2*flx12 5000p -22u*2*flx12 5001p 0 )
IINITALB11 0 INITIALB11 PWL( 0 0 20P -22u*2*flxb11 5000p -22u*2*flxb11 5001p 0)

IINITAL13 0 INITIAL13 PWL( 0 0 20P -22U*2*flx13 5000p -22U*2*flx13 5001p 0 )
IINITAL14 0 INITIAL14 PWL( 0 0 20P -22u*2*flx14 5000p 22u*2*flx14 5001p 0 )
IINITALB12 0 INITIALB12 PWL( 0 0 20P -22u*flxb12 5000p -22u*flxb12 5001p 0


##FINAL ACTIVATION - this works 

ITHRESH11 0 THRESH11 PWL(0 0 20p 23U)
#35,30,-5
ITHRESH12 0 THRESH12 PWL(0 0 20p 30U)
ITHRESH21 0 THRESH21 PWL(0 0 20p -5U)
#was like 23u
XACTfinal COMP6 A5 DOUT21 A6  DC6 DC5   DOUTFINAL1 0   DOUTFINAL2 0   DOUTFINAL3 0   DOUTFINAL4  0 DOUTFINAL5 0 DOUTFINAL6 0   THRESH21

XNEURON1 3NEURON2 INPUT11 INPUT13 INPUTB12 TARGET1 DOUTFINAL1 DOUTFINAL2 THRESH11 A3 A5 B3 B4 DC3 DC5 DCC3 DCC4  OUTPUT1 0    OUTPUT2 0 OUTPUTAXON  DELAYEDTARGETP 0  0 DELAYEDTARGETN DELAYEDTARGETP2 0   INITIAL11 INITIAL12 INITIALB11
          #x3NEURON2 INPUT1 INPUT2 INPUTBIAS TARGET DOUTFINAL1 DOUTFINAL2 THRESH XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT DCCIN DCCOUT OUTPUT OUTPUTAXON

xbfrout1 bfrsplit4 B4 DOUTFINAL3 B6 dc6 DC8  0 actfinaloutp actfinaloutn 0 0 actfinaloutp2  actfinaloutn2 0 



#xtargetdelay bfr B6 DELAYEDTARGETp b6x dc8 dc8x delayedtargetp21 0
#xtargetdelay2 bfr A6 delayedtargetp21 A6x dc8X dc8xx delayedtargetp22 0

xtargetdelay1 bfr B6 DELAYEDTARGETP b6w dc8 dc8x  delayedtargetp11 0
xtargetdelay2 bfr A6 delayedtargetp11 A6w dc8x dc8xy   0 delayedtargetp12

xtargetdelay3 bfr b6x delayedtargetp12 b6w  dc8xy dc8xxy    0 delayedtargetp13 
xtargetdelay4 bfr A6x delayedtargetp13 A6w  dc8xxy DC8Xx delayedtargetp14 0


#XDELAYin1 DELAY10 OUTPUT1 b6x b6xx A6x A6xx DC8xx DC8xxx  0 DELAYin1   DELAYin2 0
#XDELAYin1 DELAY10 OUTPUT1 b6x b6xx A6x A6xx DC8xx DC8xxx  0 DELAYin1   DELAYin2 0

XDELAYin1 DELAY163 OUTPUT1 b6x b6xx A6x A6xx DC8xx DC8xxx  0 DELAYin1   DELAYin2 0 DELAYin0 0



#XPERCEPTRON21 PERCEPTRON2LAYER2   b6xx  B7 A7 A6Xx   delayin1  actfinaloutp actfinaloutn delayedtargetp22   DC8xxx DC9 INCR21 DECR21
XPERCEPTRON21 PERCEPTRON2LAYER2   b6xx  B7 A7 A6Xx   delayin1  actfinaloutp actfinaloutn delayedtargetp14   DC8xxx DC9 INCR21 DECR21


XDELAYinb DELAY163 ADJUSTB21 B7 B7x A7 A7x DC9x DC9  0 DELAYb1 0 DELAYb2 0 DELAYb0 0
#XDELAYinb DELAY153 ADJUSTB21 B7 B7x A7 A7x DC9x DC9  0 DELAYb1 0 DELAYb2 0 DELAYb0 0


#XCONVO CONV A7 A8   DCC5 DCC4  INCR21 DECR21 SFQOUTPLUS21 SFQOUTMINUS21
XCONVO CONV A7x A8   DCC5 DCC4  INCR21 DECR21 SFQOUTPLUS21 SFQOUTMINUS21


#XPERCEPTRONb21 PERCEPTRON2LAYER2   B7  B8 A9 A8   ADJUSTB21  actfinaloutp2 actfinaloutn2 DELAYEDTARGETP2   DC9 DC10 INCRb21 DECRb21
XPERCEPTRONb21 PERCEPTRON2LAYER2   B7x  B8 A9 A8   DELAYb1  actfinaloutp2 actfinaloutn2 delayedtargetp27   DC9x DC10 INCRb21 DECRb21

XCONVb21 CONV A9 A10   DCC6 DCC5  INCRb21 DECRb21 SFQOUTPLUSb21 SFQOUTMINUSb21

XNEURON2 3NEURON2 INPUT12 INPUT14 INPUTB13 TARGET2 DOUTFINAL5 DOUTFINAL6 THRESH12 A10 A11 B8 B9 DC10 DC11 DCC6 DCC7 OUTPUT3 0  OUTPUT4 0 OUTPUTAXON2  DELAYEDTARGETP3 0  0 DELAYEDTARGETN12  DELAYEDTARGETP4  0 INITIAL13 INITIAL14 INITIALB12



#IINITAL22 0 INITIAL22 PWL( 0 0 20P flx22*2*-22.6U 5000p flx22*2*-22.6U 5001p 0 )
IINITAL22 0 INITIAL22 PWL( 0 0 20P flx22*2*-22.6U 5000p flx22*2*-22.6U )

XSTORE22 BISTORE SFQOUTPLUS22 SFQOUTMINUS22 WEIGHTL22 WEIGHTR22



#xtargetdelay3 bfr B9 DELAYEDTARGETP3 b9x dc11 dc11x delayedtargetp23 0
#xtargetdelay4 bfr A11 delayedtargetp23 A11x dc11X dc11xx delayedtargetp24 0

xtargetdelay5 bfr B9 DELAYEDTARGETP3 b9w dc11 dc11x  delayedtargetp23 0
xtargetdelay6 bfr A11 delayedtargetp23 A11w dc11x dc11Xy   0 delayedtargetp24 

xtargetdelay7 bfr b9x delayedtargetp24 b9w  dc11Xy dc11xxy    0 delayedtargetp25 
#xtargetdelay8 bfrsplit2 A11x delayedtargetp25 A11w  dc11xxy dc11Xx  delayedtargetp26 0 
xtargetdelay8 bfrsplit2 A11x delayedtargetp25 A11w  dc11xxy dc11Xx  delayedtargetp26 0 delayedtargetp27 0 


#was delay10
#XDELAYin2 DELAY14 OUTPUT3 b9x b9xx A11x A11xx DC11xx DC11xxx  0 DELAYin3   DELAYin4 0
XDELAYin2 DELAY163 OUTPUT3 b9x b9xx A11x A11xx DC11xx DC11xxx  0 DELAYin3   DELAYin4 0 DELAYin5 0


X22 SYNAPSEfastestnext2 OUTPUTAXON2 DOUT23 DOUT22  WEIGHTL22 WEIGHTR22 INITIAL22


xbfrout2 bfrsplit2 B9xx DOUTFINAL4 B10 DC11xxx DC12  0 actfinaloutp3  actfinaloutn3 0


XPERCEPTRON22 PERCEPTRON2LAYER2   B10  0 A12 A11xx   DELAYin3  actfinaloutp3 actfinaloutn3 DELAYEDTARGETP26   DC12 0 INCR22 DECR22


#ITEST 0 TESTCONV PWL (0 0 8000P 0 8002.5P 600U 8005P 0)
#xtest LSmitll_DCSFQ_PTLTX testconv SFQOUTPLUS22
XCONVO22 CONV A12 0   0 DCC7  INCR22 DECR22 SFQOUTPLUS22 SFQOUTMINUS22







.PRINT DEVII IIN1
.PRINT DEVII IIN2
#.print devii IINBIAS1


#.print devii Iactualsynbias21
#.print devii Iactualsynbias21
.print phase lstore1.x11.XNEURON1
.print phase lstore1.x12.XNEURON1
.print phase lstore1.xb11.XNEURON1
.print phase lstore1.x11.XNEURON2
.print phase lstore1.x12.XNEURON2
.print phase lstore1.xb11.XNEURON2
.print devii IINBIAS1
.PRINT PHASE LQ.XACT11.XNEURON1
.PRINT PHASE LQ.XACT11.XNEURON2




.print phase lstore1.X21
.PRINT PHASE LSTORE1.X22
.print phase lstore1.Xb21
#.print phase linput.Xb21

.PRINT PHASE LQ.X21
.PRINT PHASE LQ.X22
.PRINT PHASE LQ.Xb21

.PRINT DEVII ITARGET
.PRINT PHASE LQ.XACTfinal

#.print phase lq.xb11.XNEURON1
#.print phase lq.xb11.XNEURON2

#.print phase lq.xtargetdelay3
#.print phase lq.xtargetdelay4
#.print phase lq.xtargetdelay5
#.print phase lq.xtargetdelay6
#.print devii Iactualsynbias21
#.print phase lq.xdelay1.XDELAYinb
#.print phase lq.xdelay15.XDELAYinb


#.print phase l1_q.xincr.XPERCEPTRON21
#.print phase l2_q.xincr.XPERCEPTRON21
#.print phase l4_q.xincr.XPERCEPTRON21
#.print phase l5_q.xincr.XPERCEPTRON21
#.print phase l1_q.xincr.XPERCEPTRONb21
#.print phase l2_q.xincr.XPERCEPTRONb21
#.print phase l4_q.xincr.XPERCEPTRONb21
#.print phase l5_q.xincr.XPERCEPTRONb21
#.print phase l1_q.xdecr.XPERCEPTRONb21
#.print phase l2_q.xdecr.XPERCEPTRONb21
#.print phase l4_q.xdecr.XPERCEPTRONb21
#.print phase l5_q.xdecr.XPERCEPTRONb21



#.PRINT PHASE LQ.XACTfinal


.SUBCKT 3NEURON2 INPUT1 INPUT2 INPUTBIAS TARGET ACTNEXT1 ACTNEXT2 THRESH XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT DCCIN DCCOUT OUTPUT1 OUTPUT1GND OUTPUT2 OUTPUT2GND OUTPUTAXON DELAYOUTTARGET3 DELAYOUTTARGET3GND DELAYOUTTARGET4 DELAYOUTTARGET4GND DELAYOUTTARGET5 DELAYOUTTARGET5GND INITIAL11 INITIAL12 INITIALB11

#INPUTS
LSYN11 INPUT1 SYN11 1p  
LSYN12 INPUT2 SYN12 1p  
LSYNB11 INPUTBIAS SYNB11 1p  
LTARGET1 TARGET TARGET1 1p
LTARGET2 TARGET1 0 1p

#COUPLINGS
KSYN11 LSYN11 LSYNADJUST11 -0.1
KSYN12 LSYN12 LSYNADJUST12 -0.1
KSYNB11 LSYNB11 LSYNADJUSTB11 -0.1
KT1 LTARGET1 LADJUSTTARGET1 -0.05
KT2 LTARGET2 LADJUSTTARGET2 -0.05
LSYNADJUST11 0 ADJUST11 5P 
LSYNADJUST12 0 ADJUST12 5P 
LSYNADJUSTB11 0 ADJUSTB11 5P 
LADJUSTTARGET1 0 ADJUSTTARGET1 5P
LADJUSTTARGET2 0 ADJUSTTARGET2 5P


#SYNAPSE 1
#IINITAL11 0 INITIAL11 PWL( 0 0 20P -80U)
XSTORE11 BISTORE SFQOUTPLUS11 SFQOUTMINUS11 WEIGHTL11 WEIGHTR11
X11 SYNAPSEfastest SYN11 DOUT12 DOUT11 WEIGHTL11 WEIGHTR11 INITIAL11
#l111 SFQOUTPLUS11 0 1p
#l112 SFQOUTMINUS11 0 1p

#SYNAPSE 2
#IINITAL12 0 INITIAL12 PWL( 0 0 20P -80U)
XSTORE12 BISTORE SFQOUTPLUS12 SFQOUTMINUS12 WEIGHTL12 WEIGHTR12
X12 SYNAPSEfastest SYN12 DOUT13 DOUT12 WEIGHTL12 WEIGHTR12 INITIAL12
#l121 SFQOUTPLUS12 0 1p
#l122 SFQOUTMINUSB12 0 1p

#SYNAPSE BIAS
#IINITALB11 0 INITIALB11 PWL( 0 0 20P -80U)
XSTOREB11 BISTORE SFQOUTPLUSB11 SFQOUTMINUSB11 WEIGHTLB11 WEIGHTRB11
XB11 SYNAPSEfastest SYNB11 0 DOUT13 WEIGHTLB11 WEIGHTRB11 INITIALB11
#lB111 SFQOUTPLUSB11 0 1p
#lB112 SFQOUTMINUSB11 0 1p

#ACTIVATION
XACT11 COMP5 XIN1 DOUT11 A4 DCIN DC4 DOUTL11 0  0 DOUTR12  0 DOUTL13 OUTPUT1GND OUTPUT1 OUTPUT2GND OUTPUT2   THRESH

#AXON FOR OUTPUT
XTRANSMIT1 TRANSMIT DOUTL11 XIN2 B4 A4 A6 DC4 DC6 DCCIN DCC4 OUTPUTAXON

#DELAYS
XDELAYACT1 DELAY10 DOUTR12 B4 B5 A6 A7 DC6 DC7  DELAYOUT1 0  DELAYOUT2 0
XDELAYTARGET DELAY14 ADJUSTTARGET1 B5 B6 A7 A8 DC7 DC8  DELAYOUTTARGET1  0 DELAYOUTTARGET2 0
#XDELAYTARGET2 DELAY103 ADJUSTTARGET2 B7 B8 A9 A10 DC9 DC10  DELAYOUTTARGET3 DELAYOUTTARGET3GND   DELAYOUTTARGET4 DELAYOUTTARGET4GND DELAYOUTTARGET5  DELAYOUTTARGET5GND 
XDELAYTARGET2 DELAY143 ADJUSTTARGET2 B7 B8 A9 A10 DC9 DC10  DELAYOUTTARGET3 DELAYOUTTARGET3GND   DELAYOUTTARGET4 DELAYOUTTARGET4GND DELAYOUTTARGET5  DELAYOUTTARGET5GND 
#i think this was delay143


#LEARNING ALGORITHMS
#ASSUME DOUTFINAL1 0 DOUTFINAL2 0  DOUTFINAL3 0  0 DOUTFINAL4
#XMLP MLPNEW B6 B7 A8 A9 DELAYOUT1 DELAYOUT2 DELAYOUTTARGET1 DELAYOUTTARGET2 ACTNEXT1 ACTNEXT2 DC8 DC9 OUTPUTTARGET1L 0 OUTPUTTARGET2L 0 OUTPUTTARGET3L 0
#XDELAYTARGET2 DELAY18 ADJUSTTARGET2 B7 B8 A9 A10 DC9 dc10  DELAYOUTTARGET3GND DELAYOUTTARGET3  DELAYOUTTARGET4 DELAYOUTTARGET4GND  DELAYOUTTARGET5GND DELAYOUTTARGET5 
XMLP MLPNEW B6 B7 A8 A9 DELAYOUT1 DELAYOUT2 DELAYOUTTARGET1 DELAYOUTTARGET2 ACTNEXT1 ACTNEXT2 DC8 DC9   OUTPUTTARGET1L 0 OUTPUTTARGET2L 0 OUTPUTTARGET3L 0

XDELAYINPUT1 DELAY18 ADJUST11  B8  B9  A10 A11 DC10 DC11 DELAYOUTINPUT111 0 DELAYOUTINPUT112 0 DELAYOUTINPUT113 0 DELAYOUTINPUT114 0 DELAYOUTINPUT115 0 DELAYOUTINPUT116 0
XDELAYINPUT2 DELAY18 ADJUST12  B9  B10  A11 A12 DC11 DC12 DELAYOUTINPUT121 0 DELAYOUTINPUT122 0 DELAYOUTINPUT123 0 DELAYOUTINPUT124 0 DELAYOUTINPUT125 0 DELAYOUTINPUT126 0
XDELAYINPUTB1 DELAY18 ADJUSTB11  B10  B11  A12 A13 DC12 DC13 DELAYOUTINPUT1B1 0 DELAYOUTINPUT1B2 0 DELAYOUTINPUT1B3 0 DELAYOUTINPUT1B4 0 DELAYOUTINPUT1B5 0 DELAYOUTINPUT1B6 0

XDELAYact2 DELAY15 DOUTL13  B11 B12  A13 A14 DC13 DC14  DELAYOUTact111 0 0  DELAYOUTact112 DELAYOUTact113 0 0  DELAYOUTact114   DELAYOUTact115  0 0  DELAYOUTact116 
#XDELAYact2 DELAY15 DOUTL13  B11 B12  A13 A14 DC13 DC14  0 DELAYOUTact111 DELAYOUTact112 0 DELAYOUTact113 0 0  DELAYOUTact114   DELAYOUTact115  0 0  DELAYOUTact116 


XPERCEPTRON11 PERCEPTRON  B13 B12  A14 A15  DELAYOUTINPUT111 DELAYOUTact111 DELAYOUTact112 OUTPUTTARGET1L DC15 DC14 INCR11 DECR11
XPERCEPTRON12 PERCEPTRON  B14 B13  A15 A16  DELAYOUTINPUT121 DELAYOUTact113 DELAYOUTact114 OUTPUTTARGET2L DC16 DC15 INCR12 DECR12
XPERCEPTRONB11 PERCEPTRON  XOUT2 B14  A16 A17  DELAYOUTINPUT1B1 DELAYOUTact115 DELAYOUTact116 OUTPUTTARGET3L DCOUT DC16 INCRB11 DECRB11

XCONV11 CONV A17 A18 DCC5 DCC4 INCR11 DECR11 SFQOUTPLUS11 SFQOUTMINUS11
XCONV12 CONV A18 A19 DCC6 DCC5 INCR12 DECR12 SFQOUTPLUS12 SFQOUTMINUS12
XCONVB11 CONV A19 XOUT1 DCCOUT DCC6 INCRB11 DECRB11 SFQOUTPLUSB11 SFQOUTMINUSB11

.ENDS 3NEURON2


.SUBCKT MLPNEW XIN1 XOUT1 XIN2 XOUT2 OI1 OI2 T1 T2 OJ1 OJ2 DCIN DCOUT OUTPUTTARGET1L OUTPUTTARGET1R OUTPUTTARGET2L OUTPUTTARGET2R OUTPUTTARGET3L OUTPUTTARGET3R
#Oi.T
Xand1  AND  B7 XIN1  XIN2 A9  OI1 T1 DC9 DCIN  andout1
#Oi.!Oj
Xand2  AND B8 B7 A9 A10 OI2 OJ1 DC10 DC9 andout2
#T.!Oj
Xand3  AND B9 B8 A10 A11 T2 OJ2 DC11 DC10 andout3
#D=Oi.T + Oi.!Oj + T.!Oj 
X3OR OR3 B9 XOUT1 XOUT2 A11   ANDOUT1 ANDOUT2 ANDOUT3 DCOUT DC11  OUTPUTTARGET1L OUTPUTTARGET1R OUTPUTTARGET2L OUTPUTTARGET2R OUTPUTTARGET3L OUTPUTTARGET3R 
.ENDS MLPNEW













.SUBCKT DELAY10 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 XOUT1  DC15 DC14      DELAYOUT9 0
XDELAY10 bfrsplit2 XOUT2 DELAYOUT9 A10   DC15 DCOUT      OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R
.ends DELAY10


.SUBCKT DELAY103 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R  OUTPUT3L OUTPUT3R

XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR XOUT2 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 bfrsplit3 XOUT1 DELAYOUT6 B7  DCOUT DC12 OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R

.ends DELAY103


.SUBCKT DELAY11 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR XOUT2 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 bfrsplit2 XOUT1 DELAYOUT10 B9   DCOUT DC16   OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R

.ends DELAY11


.SUBCKT DELAY113 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR XOUT2 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 bfrsplit3 XOUT1 DELAYOUT10 B9   DCOUT DC16   OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R

.ends DELAY113




.SUBCKT DELAY14 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R

XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR A11 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 BFR B10 DELAYOUT10 B9   DC17 DC16   DELAYOUT11 0
XDELAY12 BFR A11 DELAYOUT11 A12   DC17 DC18  DELAYOUT12 0
XDELAY13 BFR B10 DELAYOUT12 XOUT1  DC19 DC18  DELAYOUT13 0
XDELAY14 bfrsplit2 XOUT2 DELAYOUT13 A12  DC19 DCOUT  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R
#XDELAY14 bfrsplit5 XOUT2 DELAYOUT13 A12  DC19 DCOUT  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R OUTPUT4L OUTPUT4R OUTPUT5L OUTPUT5R

.ends DELAY14


.SUBCKT DELAY143 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R

XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR A11 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 BFR B10 DELAYOUT10 B9   DC17 DC16   DELAYOUT11 0
XDELAY12 BFR A11 DELAYOUT11 A12   DC17 DC18  DELAYOUT12 0
XDELAY13 BFR B10 DELAYOUT12 XOUT1  DC19 DC18  DELAYOUT13 0
XDELAY14 bfrsplit3 XOUT2 DELAYOUT13 A12  DC19 DCOUT  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R
#XDELAY14 bfrsplit5 XOUT2 DELAYOUT13 A12  DC19 DCOUT  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R OUTPUT4L OUTPUT4R OUTPUT5L OUTPUT5R

.ends DELAY143

.SUBCKT DELAY15 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R OUTPUT4L OUTPUT4R OUTPUT5L OUTPUT5R OUTPUT6L OUTPUT6R
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR A11 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 BFR B10 DELAYOUT10 B9   DC17 DC16   DELAYOUT11 0
XDELAY12 BFR A11 DELAYOUT11 A12   DC17 DC18  DELAYOUT12 0
XDELAY13 BFR B10 DELAYOUT12 B11  DC19 DC18  DELAYOUT13 0
XDELAY14 BFR XOUT2 DELAYOUT13 A12  DC19 DC20  DELAYOUT14 0

XDELAY15 bfrsplit6 XOUT1 DELAYOUT14 B11 DCOUT DC20  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R OUTPUT4L OUTPUT4R OUTPUT5L OUTPUT5R OUTPUT6L OUTPUT6R

.ends DELAY15

.SUBCKT DELAY153 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R 
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR A11 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 BFR B10 DELAYOUT10 B9   DC17 DC16   DELAYOUT11 0
XDELAY12 BFR A11 DELAYOUT11 A12   DC17 DC18  DELAYOUT12 0
XDELAY13 BFR B10 DELAYOUT12 B11  DC19 DC18  DELAYOUT13 0
XDELAY14 BFR XOUT2 DELAYOUT13 A12  DC19 DC20  DELAYOUT14 0

XDELAY15 bfrsplit3 XOUT1 DELAYOUT14 B11 DCOUT DC20  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R 

.ends DELAY153



.SUBCKT DELAY16 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR A11 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 BFR B10 DELAYOUT10 B9   DC17 DC16   DELAYOUT11 0
XDELAY12 BFR A11 DELAYOUT11 A12   DC17 DC18  DELAYOUT12 0
XDELAY13 BFR B10 DELAYOUT12 B11  DC19 DC18  DELAYOUT13 0
XDELAY14 BFR A13 DELAYOUT13 A12  DC19 DC20  DELAYOUT14 0
XDELAY15 BFR XOUT1 DELAYOUT14 B11  DC21 DC20  DELAYOUT15 0
XDELAY16 bfrsplit2 A13 DELAYOUT15 XOUT2  DC21 DCOUT  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R
.ends DELAY16

.SUBCKT DELAY163 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR A11 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 BFR B10 DELAYOUT10 B9   DC17 DC16   DELAYOUT11 0
XDELAY12 BFR A11 DELAYOUT11 A12   DC17 DC18  DELAYOUT12 0
XDELAY13 BFR B10 DELAYOUT12 B11  DC19 DC18  DELAYOUT13 0
XDELAY14 BFR A13 DELAYOUT13 A12  DC19 DC20  DELAYOUT14 0
XDELAY15 BFR XOUT1 DELAYOUT14 B11  DC21 DC20  DELAYOUT15 0
XDELAY16 bfrsplit3 A13 DELAYOUT15 XOUT2  DC21 DCOUT  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R
.ends DELAY163


.SUBCKT DELAY18 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR A11 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 BFR B10 DELAYOUT10 B9   DC17 DC16   DELAYOUT11 0
XDELAY12 BFR A11 DELAYOUT11 A12   DC17 DC18  DELAYOUT12 0
XDELAY13 BFR B10 DELAYOUT12 B11  DC19 DC18  DELAYOUT13 0
XDELAY14 BFR A13 DELAYOUT13 A12  DC19 DC20  DELAYOUT14 0
XDELAY15 BFR B12 DELAYOUT14 B11  DC21 DC20  DELAYOUT15 0
XDELAY16 BFR A13 DELAYOUT15 A14  DC21 DC22  DELAYOUT16 0
XDELAY17 BFR B12 DELAYOUT16 XOUT1  DC23 DC22  DELAYOUT17 0
XDELAY18 bfrsplit3 XOUT2 DELAYOUT17 A14 DC23 DCOUT  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R  OUTPUT3L OUTPUT3R


.ends DELAY18

***    INPUTS  ***
IIN1 0 IN1 PWL(0 0 20P 0 1.55000e-09 0.00000e+00 1.55500e-09 2.00000e-03 1.60500e-09 2.00000e-03
+ 1.61000e-09 0.00000e+00 3.55000e-09 0.00000e+00 3.55500e-09 2.00000e-03
+ 3.60500e-09 2.00000e-03 3.61000e-09 0.00000e+00 5.55000e-09 0.00000e+00
+ 5.55500e-09 2.00000e-03 5.60500e-09 2.00000e-03 5.61000e-09 0.00000e+00
+ 7.55000e-09 0.00000e+00 7.55500e-09 2.00000e-03 7.60500e-09 2.00000e-03
+ 7.61000e-09 0.00000e+00 9.55000e-09 0.00000e+00 9.55500e-09 2.00000e-03
+ 9.60500e-09 2.00000e-03 9.61000e-09 0.00000e+00 1.15500e-08 0.00000e+00
+ 1.15550e-08 2.00000e-03 1.16050e-08 2.00000e-03 1.16100e-08 0.00000e+00
+ 1.35500e-08 0.00000e+00 1.35550e-08 2.00000e-03 1.36050e-08 2.00000e-03
+ 1.36100e-08 0.00000e+00 1.55500e-08 0.00000e+00 1.55550e-08 2.00000e-03
+ 1.56050e-08 2.00000e-03 1.56100e-08 0.00000e+00 1.75500e-08 0.00000e+00
+ 1.75550e-08 2.00000e-03 1.76050e-08 2.00000e-03 1.76100e-08 0.00000e+00
+ 1.95500e-08 0.00000e+00 1.95550e-08 2.00000e-03 1.96050e-08 2.00000e-03
+ 1.96100e-08 0.00000e+00 2.15500e-08 0.00000e+00 2.15550e-08 2.00000e-03
+ 2.16050e-08 2.00000e-03 2.16100e-08 0.00000e+00 2.35500e-08 0.00000e+00
+ 2.35550e-08 2.00000e-03 2.36050e-08 2.00000e-03 2.36100e-08 0.00000e+00
+ 2.55500e-08 0.00000e+00 2.55550e-08 2.00000e-03 2.56050e-08 2.00000e-03
+ 2.56100e-08 0.00000e+00 2.75500e-08 0.00000e+00 2.75550e-08 2.00000e-03
+ 2.76050e-08 2.00000e-03 2.76100e-08 0.00000e+00 2.95500e-08 0.00000e+00
+ 2.95550e-08 2.00000e-03 2.96050e-08 2.00000e-03 2.96100e-08 0.00000e+00
+ 3.15500e-08 0.00000e+00 3.15550e-08 2.00000e-03 3.16050e-08 2.00000e-03
+ 3.16100e-08 0.00000e+00 3.35500e-08 0.00000e+00 3.35550e-08 2.00000e-03
+ 3.36050e-08 2.00000e-03 3.36100e-08 0.00000e+00 3.55500e-08 0.00000e+00
+ 3.55550e-08 2.00000e-03 3.56050e-08 2.00000e-03 3.56100e-08 0.00000e+00
+ 3.75500e-08 0.00000e+00 3.75550e-08 2.00000e-03 3.76050e-08 2.00000e-03
+ 3.76100e-08 0.00000e+00 3.95500e-08 0.00000e+00 3.95550e-08 2.00000e-03
+ 3.96050e-08 2.00000e-03 3.96100e-08 0.00000e+00 4.15500e-08 0.00000e+00
+ 4.15550e-08 2.00000e-03 4.16050e-08 2.00000e-03 4.16100e-08 0.00000e+00
+ 4.35500e-08 0.00000e+00 4.35550e-08 2.00000e-03 4.36050e-08 2.00000e-03
+ 4.36100e-08 0.00000e+00 4.55500e-08 0.00000e+00 4.55550e-08 2.00000e-03
+ 4.56050e-08 2.00000e-03 4.56100e-08 0.00000e+00 4.75500e-08 0.00000e+00
+ 4.75550e-08 2.00000e-03 4.76050e-08 2.00000e-03 4.76100e-08 0.00000e+00
+ 4.95500e-08 0.00000e+00 4.95550e-08 2.00000e-03 4.96050e-08 2.00000e-03
+ 4.96100e-08 0.00000e+00 5.15500e-08 0.00000e+00 5.15550e-08 2.00000e-03
+ 5.16050e-08 2.00000e-03 5.16100e-08 0.00000e+00 5.35500e-08 0.00000e+00
+ 5.35550e-08 2.00000e-03 5.36050e-08 2.00000e-03 5.36100e-08 0.00000e+00
+ 5.55500e-08 0.00000e+00 5.55550e-08 2.00000e-03 5.56050e-08 2.00000e-03
+ 5.56100e-08 0.00000e+00 5.75500e-08 0.00000e+00 5.75550e-08 2.00000e-03
+ 5.76050e-08 2.00000e-03 5.76100e-08 0.00000e+00 5.95500e-08 0.00000e+00
+ 5.95550e-08 2.00000e-03 5.96050e-08 2.00000e-03 5.96100e-08 0.00000e+00
+ 6.15500e-08 0.00000e+00 6.15550e-08 2.00000e-03 6.16050e-08 2.00000e-03
+ 6.16100e-08 0.00000e+00 6.35500e-08 0.00000e+00 6.35550e-08 2.00000e-03
+ 6.36050e-08 2.00000e-03 6.36100e-08 0.00000e+00 6.55500e-08 0.00000e+00
+ 6.55550e-08 2.00000e-03 6.56050e-08 2.00000e-03 6.56100e-08 0.00000e+00
+ 6.75500e-08 0.00000e+00 6.75550e-08 2.00000e-03 6.76050e-08 2.00000e-03
+ 6.76100e-08 0.00000e+00 6.95500e-08 0.00000e+00 6.95550e-08 2.00000e-03
+ 6.96050e-08 2.00000e-03 6.96100e-08 0.00000e+00 7.15500e-08 0.00000e+00
+ 7.15550e-08 2.00000e-03 7.16050e-08 2.00000e-03 7.16100e-08 0.00000e+00
+ 7.35500e-08 0.00000e+00 7.35550e-08 2.00000e-03 7.36050e-08 2.00000e-03
+ 7.36100e-08 0.00000e+00 7.55500e-08 0.00000e+00 7.55550e-08 2.00000e-03
+ 7.56050e-08 2.00000e-03 7.56100e-08 0.00000e+00 7.75500e-08 0.00000e+00
+ 7.75550e-08 2.00000e-03 7.76050e-08 2.00000e-03 7.76100e-08 0.00000e+00
+ 7.95500e-08 0.00000e+00 7.95550e-08 2.00000e-03 7.96050e-08 2.00000e-03
+ 7.96100e-08 0.00000e+00 8.15500e-08 0.00000e+00 8.15550e-08 2.00000e-03
+ 8.16050e-08 2.00000e-03 8.16100e-08 0.00000e+00 8.35500e-08 0.00000e+00
+ 8.35550e-08 2.00000e-03 8.36050e-08 2.00000e-03 8.36100e-08 0.00000e+00
+ 8.55500e-08 0.00000e+00 8.55550e-08 2.00000e-03 8.56050e-08 2.00000e-03
+ 8.56100e-08 0.00000e+00 8.75500e-08 0.00000e+00 8.75550e-08 2.00000e-03
+ 8.76050e-08 2.00000e-03 8.76100e-08 0.00000e+00 8.95500e-08 0.00000e+00
+ 8.95550e-08 2.00000e-03 8.96050e-08 2.00000e-03 8.96100e-08 0.00000e+00
+ 9.15500e-08 0.00000e+00 9.15550e-08 2.00000e-03 9.16050e-08 2.00000e-03
+ 9.16100e-08 0.00000e+00 9.35500e-08 0.00000e+00 9.35550e-08 2.00000e-03
+ 9.36050e-08 2.00000e-03 9.36100e-08 0.00000e+00 9.55500e-08 0.00000e+00
+ 9.55550e-08 2.00000e-03 9.56050e-08 2.00000e-03 9.56100e-08 0.00000e+00
+ 9.75500e-08 0.00000e+00 9.75550e-08 2.00000e-03 9.76050e-08 2.00000e-03
+ 9.76100e-08 0.00000e+00 9.95500e-08 0.00000e+00 9.95550e-08 2.00000e-03
+ 9.96050e-08 2.00000e-03 9.96100e-08 0.00000e+00 1.01550e-07 0.00000e+00
+ 1.01555e-07 2.00000e-03 1.01605e-07 2.00000e-03 1.01610e-07 0.00000e+00
+ 1.03550e-07 0.00000e+00 1.03555e-07 2.00000e-03 1.03605e-07 2.00000e-03
+ 1.03610e-07 0.00000e+00 1.05550e-07 0.00000e+00 1.05555e-07 2.00000e-03
+ 1.05605e-07 2.00000e-03 1.05610e-07 0.00000e+00 1.07550e-07 0.00000e+00
+ 1.07555e-07 2.00000e-03 1.07605e-07 2.00000e-03 1.07610e-07 0.00000e+00
+ 1.09550e-07 0.00000e+00 1.09555e-07 2.00000e-03 1.09605e-07 2.00000e-03
+ 1.09610e-07 0.00000e+00 1.11550e-07 0.00000e+00 1.11555e-07 2.00000e-03
+ 1.11605e-07 2.00000e-03 1.11610e-07 0.00000e+00 1.13550e-07 0.00000e+00
+ 1.13555e-07 2.00000e-03 1.13605e-07 2.00000e-03 1.13610e-07 0.00000e+00
+ 1.15550e-07 0.00000e+00 1.15555e-07 2.00000e-03 1.15605e-07 2.00000e-03
+ 1.15610e-07 0.00000e+00 1.17550e-07 0.00000e+00 1.17555e-07 2.00000e-03
+ 1.17605e-07 2.00000e-03 1.17610e-07 0.00000e+00 1.19550e-07 0.00000e+00
+ 1.19555e-07 2.00000e-03 1.19605e-07 2.00000e-03 1.19610e-07 0.00000e+00
+ 1.21550e-07 0.00000e+00 1.21555e-07 2.00000e-03 1.21605e-07 2.00000e-03
+ 1.21610e-07 0.00000e+00 1.23550e-07 0.00000e+00 1.23555e-07 2.00000e-03
+ 1.23605e-07 2.00000e-03 1.23610e-07 0.00000e+00 1.25550e-07 0.00000e+00
+ 1.25555e-07 2.00000e-03 1.25605e-07 2.00000e-03 1.25610e-07 0.00000e+00
+ 1.27550e-07 0.00000e+00 1.27555e-07 2.00000e-03 1.27605e-07 2.00000e-03
+ 1.27610e-07 0.00000e+00 1.29550e-07 0.00000e+00 1.29555e-07 2.00000e-03
+ 1.29605e-07 2.00000e-03 1.29610e-07 0.00000e+00 1.31550e-07 0.00000e+00
+ 1.31555e-07 2.00000e-03 1.31605e-07 2.00000e-03 1.31610e-07 0.00000e+00
+ 1.33550e-07 0.00000e+00 1.33555e-07 2.00000e-03 1.33605e-07 2.00000e-03
+ 1.33610e-07 0.00000e+00 1.35550e-07 0.00000e+00 1.35555e-07 2.00000e-03
+ 1.35605e-07 2.00000e-03 1.35610e-07 0.00000e+00 1.37550e-07 0.00000e+00
+ 1.37555e-07 2.00000e-03 1.37605e-07 2.00000e-03 1.37610e-07 0.00000e+00
+ 1.39550e-07 0.00000e+00 1.39555e-07 2.00000e-03 1.39605e-07 2.00000e-03
+ 1.39610e-07 0.00000e+00 1.41550e-07 0.00000e+00 1.41555e-07 2.00000e-03
+ 1.41605e-07 2.00000e-03 1.41610e-07 0.00000e+00 1.43550e-07 0.00000e+00
+ 1.43555e-07 2.00000e-03 1.43605e-07 2.00000e-03 1.43610e-07 0.00000e+00
+ 1.45550e-07 0.00000e+00 1.45555e-07 2.00000e-03 1.45605e-07 2.00000e-03
+ 1.45610e-07 0.00000e+00 1.47550e-07 0.00000e+00 1.47555e-07 2.00000e-03
+ 1.47605e-07 2.00000e-03 1.47610e-07 0.00000e+00 1.49550e-07 0.00000e+00
+ 1.49555e-07 2.00000e-03 1.49605e-07 2.00000e-03 1.49610e-07 0.00000e+00
+ 1.51550e-07 0.00000e+00 1.51555e-07 2.00000e-03 1.51605e-07 2.00000e-03
+ 1.51610e-07 0.00000e+00 1.53550e-07 0.00000e+00 1.53555e-07 2.00000e-03
+ 1.53605e-07 2.00000e-03 1.53610e-07 0.00000e+00 1.55550e-07 0.00000e+00
+ 1.55555e-07 2.00000e-03 1.55605e-07 2.00000e-03 1.55610e-07 0.00000e+00
+ 1.57550e-07 0.00000e+00 1.57555e-07 2.00000e-03 1.57605e-07 2.00000e-03
+ 1.57610e-07 0.00000e+00 1.59550e-07 0.00000e+00 1.59555e-07 2.00000e-03
+ 1.59605e-07 2.00000e-03 1.59610e-07 0.00000e+00 1.61550e-07 0.00000e+00
+ 1.61555e-07 2.00000e-03 1.61605e-07 2.00000e-03 1.61610e-07 0.00000e+00
+ 1.63550e-07 0.00000e+00 1.63555e-07 2.00000e-03 1.63605e-07 2.00000e-03
+ 1.63610e-07 0.00000e+00 1.65550e-07 0.00000e+00 1.65555e-07 2.00000e-03
+ 1.65605e-07 2.00000e-03 1.65610e-07 0.00000e+00 1.67550e-07 0.00000e+00
+ 1.67555e-07 2.00000e-03 1.67605e-07 2.00000e-03 1.67610e-07 0.00000e+00
+ 1.69550e-07 0.00000e+00 1.69555e-07 2.00000e-03 1.69605e-07 2.00000e-03
+ 1.69610e-07 0.00000e+00 1.71550e-07 0.00000e+00 1.71555e-07 2.00000e-03
+ 1.71605e-07 2.00000e-03 1.71610e-07 0.00000e+00 1.73550e-07 0.00000e+00
+ 1.73555e-07 2.00000e-03 1.73605e-07 2.00000e-03 1.73610e-07 0.00000e+00
+ 1.75550e-07 0.00000e+00 1.75555e-07 2.00000e-03 1.75605e-07 2.00000e-03
+ 1.75610e-07 0.00000e+00 1.77550e-07 0.00000e+00 1.77555e-07 2.00000e-03
+ 1.77605e-07 2.00000e-03 1.77610e-07 0.00000e+00 1.79550e-07 0.00000e+00
+ 1.79555e-07 2.00000e-03 1.79605e-07 2.00000e-03 1.79610e-07 0.00000e+00
+ 1.81550e-07 0.00000e+00 1.81555e-07 2.00000e-03 1.81605e-07 2.00000e-03
+ 1.81610e-07 0.00000e+00 1.83550e-07 0.00000e+00 1.83555e-07 2.00000e-03
+ 1.83605e-07 2.00000e-03 1.83610e-07 0.00000e+00 1.85550e-07 0.00000e+00
+ 1.85555e-07 2.00000e-03 1.85605e-07 2.00000e-03 1.85610e-07 0.00000e+00
+ 1.87550e-07 0.00000e+00 1.87555e-07 2.00000e-03 1.87605e-07 2.00000e-03
+ 1.87610e-07 0.00000e+00 1.89550e-07 0.00000e+00 1.89555e-07 2.00000e-03
+ 1.89605e-07 2.00000e-03 1.89610e-07 0.00000e+00 1.91550e-07 0.00000e+00
+ 1.91555e-07 2.00000e-03 1.91605e-07 2.00000e-03 1.91610e-07 0.00000e+00
+ 1.93550e-07 0.00000e+00 1.93555e-07 2.00000e-03 1.93605e-07 2.00000e-03
+ 1.93610e-07 0.00000e+00 1.95550e-07 0.00000e+00 1.95555e-07 2.00000e-03
+ 1.95605e-07 2.00000e-03 1.95610e-07 0.00000e+00 1.97550e-07 0.00000e+00
+ 1.97555e-07 2.00000e-03 1.97605e-07 2.00000e-03 1.97610e-07 0.00000e+00
+ 1.99550e-07 0.00000e+00 1.99555e-07 2.00000e-03 1.99605e-07 2.00000e-03
+ 1.99610e-07 0.00000e+00)
IIN2 0 IN2 PWL(0 0 20P 0 2.55000e-09 0.00000e+00 2.55500e-09 2.00000e-03 2.60500e-09 2.00000e-03
+ 2.61000e-09 0.00000e+00 3.55000e-09 0.00000e+00 3.55500e-09 2.00000e-03
+ 3.60500e-09 2.00000e-03 3.61000e-09 0.00000e+00 6.55000e-09 0.00000e+00
+ 6.55500e-09 2.00000e-03 6.60500e-09 2.00000e-03 6.61000e-09 0.00000e+00
+ 7.55000e-09 0.00000e+00 7.55500e-09 2.00000e-03 7.60500e-09 2.00000e-03
+ 7.61000e-09 0.00000e+00 1.05500e-08 0.00000e+00 1.05550e-08 2.00000e-03
+ 1.06050e-08 2.00000e-03 1.06100e-08 0.00000e+00 1.15500e-08 0.00000e+00
+ 1.15550e-08 2.00000e-03 1.16050e-08 2.00000e-03 1.16100e-08 0.00000e+00
+ 1.45500e-08 0.00000e+00 1.45550e-08 2.00000e-03 1.46050e-08 2.00000e-03
+ 1.46100e-08 0.00000e+00 1.55500e-08 0.00000e+00 1.55550e-08 2.00000e-03
+ 1.56050e-08 2.00000e-03 1.56100e-08 0.00000e+00 1.85500e-08 0.00000e+00
+ 1.85550e-08 2.00000e-03 1.86050e-08 2.00000e-03 1.86100e-08 0.00000e+00
+ 1.95500e-08 0.00000e+00 1.95550e-08 2.00000e-03 1.96050e-08 2.00000e-03
+ 1.96100e-08 0.00000e+00 2.25500e-08 0.00000e+00 2.25550e-08 2.00000e-03
+ 2.26050e-08 2.00000e-03 2.26100e-08 0.00000e+00 2.35500e-08 0.00000e+00
+ 2.35550e-08 2.00000e-03 2.36050e-08 2.00000e-03 2.36100e-08 0.00000e+00
+ 2.65500e-08 0.00000e+00 2.65550e-08 2.00000e-03 2.66050e-08 2.00000e-03
+ 2.66100e-08 0.00000e+00 2.75500e-08 0.00000e+00 2.75550e-08 2.00000e-03
+ 2.76050e-08 2.00000e-03 2.76100e-08 0.00000e+00 3.05500e-08 0.00000e+00
+ 3.05550e-08 2.00000e-03 3.06050e-08 2.00000e-03 3.06100e-08 0.00000e+00
+ 3.15500e-08 0.00000e+00 3.15550e-08 2.00000e-03 3.16050e-08 2.00000e-03
+ 3.16100e-08 0.00000e+00 3.45500e-08 0.00000e+00 3.45550e-08 2.00000e-03
+ 3.46050e-08 2.00000e-03 3.46100e-08 0.00000e+00 3.55500e-08 0.00000e+00
+ 3.55550e-08 2.00000e-03 3.56050e-08 2.00000e-03 3.56100e-08 0.00000e+00
+ 3.85500e-08 0.00000e+00 3.85550e-08 2.00000e-03 3.86050e-08 2.00000e-03
+ 3.86100e-08 0.00000e+00 3.95500e-08 0.00000e+00 3.95550e-08 2.00000e-03
+ 3.96050e-08 2.00000e-03 3.96100e-08 0.00000e+00 4.25500e-08 0.00000e+00
+ 4.25550e-08 2.00000e-03 4.26050e-08 2.00000e-03 4.26100e-08 0.00000e+00
+ 4.35500e-08 0.00000e+00 4.35550e-08 2.00000e-03 4.36050e-08 2.00000e-03
+ 4.36100e-08 0.00000e+00 4.65500e-08 0.00000e+00 4.65550e-08 2.00000e-03
+ 4.66050e-08 2.00000e-03 4.66100e-08 0.00000e+00 4.75500e-08 0.00000e+00
+ 4.75550e-08 2.00000e-03 4.76050e-08 2.00000e-03 4.76100e-08 0.00000e+00
+ 5.05500e-08 0.00000e+00 5.05550e-08 2.00000e-03 5.06050e-08 2.00000e-03
+ 5.06100e-08 0.00000e+00 5.15500e-08 0.00000e+00 5.15550e-08 2.00000e-03
+ 5.16050e-08 2.00000e-03 5.16100e-08 0.00000e+00 5.45500e-08 0.00000e+00
+ 5.45550e-08 2.00000e-03 5.46050e-08 2.00000e-03 5.46100e-08 0.00000e+00
+ 5.55500e-08 0.00000e+00 5.55550e-08 2.00000e-03 5.56050e-08 2.00000e-03
+ 5.56100e-08 0.00000e+00 5.85500e-08 0.00000e+00 5.85550e-08 2.00000e-03
+ 5.86050e-08 2.00000e-03 5.86100e-08 0.00000e+00 5.95500e-08 0.00000e+00
+ 5.95550e-08 2.00000e-03 5.96050e-08 2.00000e-03 5.96100e-08 0.00000e+00
+ 6.25500e-08 0.00000e+00 6.25550e-08 2.00000e-03 6.26050e-08 2.00000e-03
+ 6.26100e-08 0.00000e+00 6.35500e-08 0.00000e+00 6.35550e-08 2.00000e-03
+ 6.36050e-08 2.00000e-03 6.36100e-08 0.00000e+00 6.65500e-08 0.00000e+00
+ 6.65550e-08 2.00000e-03 6.66050e-08 2.00000e-03 6.66100e-08 0.00000e+00
+ 6.75500e-08 0.00000e+00 6.75550e-08 2.00000e-03 6.76050e-08 2.00000e-03
+ 6.76100e-08 0.00000e+00 7.05500e-08 0.00000e+00 7.05550e-08 2.00000e-03
+ 7.06050e-08 2.00000e-03 7.06100e-08 0.00000e+00 7.15500e-08 0.00000e+00
+ 7.15550e-08 2.00000e-03 7.16050e-08 2.00000e-03 7.16100e-08 0.00000e+00
+ 7.45500e-08 0.00000e+00 7.45550e-08 2.00000e-03 7.46050e-08 2.00000e-03
+ 7.46100e-08 0.00000e+00 7.55500e-08 0.00000e+00 7.55550e-08 2.00000e-03
+ 7.56050e-08 2.00000e-03 7.56100e-08 0.00000e+00 7.85500e-08 0.00000e+00
+ 7.85550e-08 2.00000e-03 7.86050e-08 2.00000e-03 7.86100e-08 0.00000e+00
+ 7.95500e-08 0.00000e+00 7.95550e-08 2.00000e-03 7.96050e-08 2.00000e-03
+ 7.96100e-08 0.00000e+00 8.25500e-08 0.00000e+00 8.25550e-08 2.00000e-03
+ 8.26050e-08 2.00000e-03 8.26100e-08 0.00000e+00 8.35500e-08 0.00000e+00
+ 8.35550e-08 2.00000e-03 8.36050e-08 2.00000e-03 8.36100e-08 0.00000e+00
+ 8.65500e-08 0.00000e+00 8.65550e-08 2.00000e-03 8.66050e-08 2.00000e-03
+ 8.66100e-08 0.00000e+00 8.75500e-08 0.00000e+00 8.75550e-08 2.00000e-03
+ 8.76050e-08 2.00000e-03 8.76100e-08 0.00000e+00 9.05500e-08 0.00000e+00
+ 9.05550e-08 2.00000e-03 9.06050e-08 2.00000e-03 9.06100e-08 0.00000e+00
+ 9.15500e-08 0.00000e+00 9.15550e-08 2.00000e-03 9.16050e-08 2.00000e-03
+ 9.16100e-08 0.00000e+00 9.45500e-08 0.00000e+00 9.45550e-08 2.00000e-03
+ 9.46050e-08 2.00000e-03 9.46100e-08 0.00000e+00 9.55500e-08 0.00000e+00
+ 9.55550e-08 2.00000e-03 9.56050e-08 2.00000e-03 9.56100e-08 0.00000e+00
+ 9.85500e-08 0.00000e+00 9.85550e-08 2.00000e-03 9.86050e-08 2.00000e-03
+ 9.86100e-08 0.00000e+00 9.95500e-08 0.00000e+00 9.95550e-08 2.00000e-03
+ 9.96050e-08 2.00000e-03 9.96100e-08 0.00000e+00 1.02550e-07 0.00000e+00
+ 1.02555e-07 2.00000e-03 1.02605e-07 2.00000e-03 1.02610e-07 0.00000e+00
+ 1.03550e-07 0.00000e+00 1.03555e-07 2.00000e-03 1.03605e-07 2.00000e-03
+ 1.03610e-07 0.00000e+00 1.06550e-07 0.00000e+00 1.06555e-07 2.00000e-03
+ 1.06605e-07 2.00000e-03 1.06610e-07 0.00000e+00 1.07550e-07 0.00000e+00
+ 1.07555e-07 2.00000e-03 1.07605e-07 2.00000e-03 1.07610e-07 0.00000e+00
+ 1.10550e-07 0.00000e+00 1.10555e-07 2.00000e-03 1.10605e-07 2.00000e-03
+ 1.10610e-07 0.00000e+00 1.11550e-07 0.00000e+00 1.11555e-07 2.00000e-03
+ 1.11605e-07 2.00000e-03 1.11610e-07 0.00000e+00 1.14550e-07 0.00000e+00
+ 1.14555e-07 2.00000e-03 1.14605e-07 2.00000e-03 1.14610e-07 0.00000e+00
+ 1.15550e-07 0.00000e+00 1.15555e-07 2.00000e-03 1.15605e-07 2.00000e-03
+ 1.15610e-07 0.00000e+00 1.18550e-07 0.00000e+00 1.18555e-07 2.00000e-03
+ 1.18605e-07 2.00000e-03 1.18610e-07 0.00000e+00 1.19550e-07 0.00000e+00
+ 1.19555e-07 2.00000e-03 1.19605e-07 2.00000e-03 1.19610e-07 0.00000e+00
+ 1.22550e-07 0.00000e+00 1.22555e-07 2.00000e-03 1.22605e-07 2.00000e-03
+ 1.22610e-07 0.00000e+00 1.23550e-07 0.00000e+00 1.23555e-07 2.00000e-03
+ 1.23605e-07 2.00000e-03 1.23610e-07 0.00000e+00 1.26550e-07 0.00000e+00
+ 1.26555e-07 2.00000e-03 1.26605e-07 2.00000e-03 1.26610e-07 0.00000e+00
+ 1.27550e-07 0.00000e+00 1.27555e-07 2.00000e-03 1.27605e-07 2.00000e-03
+ 1.27610e-07 0.00000e+00 1.30550e-07 0.00000e+00 1.30555e-07 2.00000e-03
+ 1.30605e-07 2.00000e-03 1.30610e-07 0.00000e+00 1.31550e-07 0.00000e+00
+ 1.31555e-07 2.00000e-03 1.31605e-07 2.00000e-03 1.31610e-07 0.00000e+00
+ 1.34550e-07 0.00000e+00 1.34555e-07 2.00000e-03 1.34605e-07 2.00000e-03
+ 1.34610e-07 0.00000e+00 1.35550e-07 0.00000e+00 1.35555e-07 2.00000e-03
+ 1.35605e-07 2.00000e-03 1.35610e-07 0.00000e+00 1.38550e-07 0.00000e+00
+ 1.38555e-07 2.00000e-03 1.38605e-07 2.00000e-03 1.38610e-07 0.00000e+00
+ 1.39550e-07 0.00000e+00 1.39555e-07 2.00000e-03 1.39605e-07 2.00000e-03
+ 1.39610e-07 0.00000e+00 1.42550e-07 0.00000e+00 1.42555e-07 2.00000e-03
+ 1.42605e-07 2.00000e-03 1.42610e-07 0.00000e+00 1.43550e-07 0.00000e+00
+ 1.43555e-07 2.00000e-03 1.43605e-07 2.00000e-03 1.43610e-07 0.00000e+00
+ 1.46550e-07 0.00000e+00 1.46555e-07 2.00000e-03 1.46605e-07 2.00000e-03
+ 1.46610e-07 0.00000e+00 1.47550e-07 0.00000e+00 1.47555e-07 2.00000e-03
+ 1.47605e-07 2.00000e-03 1.47610e-07 0.00000e+00 1.50550e-07 0.00000e+00
+ 1.50555e-07 2.00000e-03 1.50605e-07 2.00000e-03 1.50610e-07 0.00000e+00
+ 1.51550e-07 0.00000e+00 1.51555e-07 2.00000e-03 1.51605e-07 2.00000e-03
+ 1.51610e-07 0.00000e+00 1.54550e-07 0.00000e+00 1.54555e-07 2.00000e-03
+ 1.54605e-07 2.00000e-03 1.54610e-07 0.00000e+00 1.55550e-07 0.00000e+00
+ 1.55555e-07 2.00000e-03 1.55605e-07 2.00000e-03 1.55610e-07 0.00000e+00
+ 1.58550e-07 0.00000e+00 1.58555e-07 2.00000e-03 1.58605e-07 2.00000e-03
+ 1.58610e-07 0.00000e+00 1.59550e-07 0.00000e+00 1.59555e-07 2.00000e-03
+ 1.59605e-07 2.00000e-03 1.59610e-07 0.00000e+00 1.62550e-07 0.00000e+00
+ 1.62555e-07 2.00000e-03 1.62605e-07 2.00000e-03 1.62610e-07 0.00000e+00
+ 1.63550e-07 0.00000e+00 1.63555e-07 2.00000e-03 1.63605e-07 2.00000e-03
+ 1.63610e-07 0.00000e+00 1.66550e-07 0.00000e+00 1.66555e-07 2.00000e-03
+ 1.66605e-07 2.00000e-03 1.66610e-07 0.00000e+00 1.67550e-07 0.00000e+00
+ 1.67555e-07 2.00000e-03 1.67605e-07 2.00000e-03 1.67610e-07 0.00000e+00
+ 1.70550e-07 0.00000e+00 1.70555e-07 2.00000e-03 1.70605e-07 2.00000e-03
+ 1.70610e-07 0.00000e+00 1.71550e-07 0.00000e+00 1.71555e-07 2.00000e-03
+ 1.71605e-07 2.00000e-03 1.71610e-07 0.00000e+00 1.74550e-07 0.00000e+00
+ 1.74555e-07 2.00000e-03 1.74605e-07 2.00000e-03 1.74610e-07 0.00000e+00
+ 1.75550e-07 0.00000e+00 1.75555e-07 2.00000e-03 1.75605e-07 2.00000e-03
+ 1.75610e-07 0.00000e+00 1.78550e-07 0.00000e+00 1.78555e-07 2.00000e-03
+ 1.78605e-07 2.00000e-03 1.78610e-07 0.00000e+00 1.79550e-07 0.00000e+00
+ 1.79555e-07 2.00000e-03 1.79605e-07 2.00000e-03 1.79610e-07 0.00000e+00
+ 1.82550e-07 0.00000e+00 1.82555e-07 2.00000e-03 1.82605e-07 2.00000e-03
+ 1.82610e-07 0.00000e+00 1.83550e-07 0.00000e+00 1.83555e-07 2.00000e-03
+ 1.83605e-07 2.00000e-03 1.83610e-07 0.00000e+00 1.86550e-07 0.00000e+00
+ 1.86555e-07 2.00000e-03 1.86605e-07 2.00000e-03 1.86610e-07 0.00000e+00
+ 1.87550e-07 0.00000e+00 1.87555e-07 2.00000e-03 1.87605e-07 2.00000e-03
+ 1.87610e-07 0.00000e+00 1.90550e-07 0.00000e+00 1.90555e-07 2.00000e-03
+ 1.90605e-07 2.00000e-03 1.90610e-07 0.00000e+00 1.91550e-07 0.00000e+00
+ 1.91555e-07 2.00000e-03 1.91605e-07 2.00000e-03 1.91610e-07 0.00000e+00
+ 1.94550e-07 0.00000e+00 1.94555e-07 2.00000e-03 1.94605e-07 2.00000e-03
+ 1.94610e-07 0.00000e+00 1.95550e-07 0.00000e+00 1.95555e-07 2.00000e-03
+ 1.95605e-07 2.00000e-03 1.95610e-07 0.00000e+00 1.98550e-07 0.00000e+00
+ 1.98555e-07 2.00000e-03 1.98605e-07 2.00000e-03 1.98610e-07 0.00000e+00
+ 1.99550e-07 0.00000e+00 1.99555e-07 2.00000e-03 1.99605e-07 2.00000e-03
+ 1.99610e-07 0.00000e+00)
IINBIAS1 0 INB11 pulse(0 0.002 550p 5p 5p 50p 1000p)
ITARGET 0 TARGET0  PWL(0 0 20P 0 5.50000e-10 0.00000e+00 5.55000e-10 2.00000e-03 6.05000e-10 2.00000e-03
+ 6.10000e-10 0.00000e+00 3.55000e-09 0.00000e+00 3.55500e-09 2.00000e-03
+ 3.60500e-09 2.00000e-03 3.61000e-09 0.00000e+00 4.55000e-09 0.00000e+00
+ 4.55500e-09 2.00000e-03 4.60500e-09 2.00000e-03 4.61000e-09 0.00000e+00
+ 7.55000e-09 0.00000e+00 7.55500e-09 2.00000e-03 7.60500e-09 2.00000e-03
+ 7.61000e-09 0.00000e+00 8.55000e-09 0.00000e+00 8.55500e-09 2.00000e-03
+ 8.60500e-09 2.00000e-03 8.61000e-09 0.00000e+00 1.15500e-08 0.00000e+00
+ 1.15550e-08 2.00000e-03 1.16050e-08 2.00000e-03 1.16100e-08 0.00000e+00
+ 1.25500e-08 0.00000e+00 1.25550e-08 2.00000e-03 1.26050e-08 2.00000e-03
+ 1.26100e-08 0.00000e+00 1.55500e-08 0.00000e+00 1.55550e-08 2.00000e-03
+ 1.56050e-08 2.00000e-03 1.56100e-08 0.00000e+00 1.65500e-08 0.00000e+00
+ 1.65550e-08 2.00000e-03 1.66050e-08 2.00000e-03 1.66100e-08 0.00000e+00
+ 1.95500e-08 0.00000e+00 1.95550e-08 2.00000e-03 1.96050e-08 2.00000e-03
+ 1.96100e-08 0.00000e+00 2.05500e-08 0.00000e+00 2.05550e-08 2.00000e-03
+ 2.06050e-08 2.00000e-03 2.06100e-08 0.00000e+00 2.35500e-08 0.00000e+00
+ 2.35550e-08 2.00000e-03 2.36050e-08 2.00000e-03 2.36100e-08 0.00000e+00
+ 2.45500e-08 0.00000e+00 2.45550e-08 2.00000e-03 2.46050e-08 2.00000e-03
+ 2.46100e-08 0.00000e+00 2.75500e-08 0.00000e+00 2.75550e-08 2.00000e-03
+ 2.76050e-08 2.00000e-03 2.76100e-08 0.00000e+00 2.85500e-08 0.00000e+00
+ 2.85550e-08 2.00000e-03 2.86050e-08 2.00000e-03 2.86100e-08 0.00000e+00
+ 3.15500e-08 0.00000e+00 3.15550e-08 2.00000e-03 3.16050e-08 2.00000e-03
+ 3.16100e-08 0.00000e+00 3.25500e-08 0.00000e+00 3.25550e-08 2.00000e-03
+ 3.26050e-08 2.00000e-03 3.26100e-08 0.00000e+00 3.55500e-08 0.00000e+00
+ 3.55550e-08 2.00000e-03 3.56050e-08 2.00000e-03 3.56100e-08 0.00000e+00
+ 3.65500e-08 0.00000e+00 3.65550e-08 2.00000e-03 3.66050e-08 2.00000e-03
+ 3.66100e-08 0.00000e+00 3.95500e-08 0.00000e+00 3.95550e-08 2.00000e-03
+ 3.96050e-08 2.00000e-03 3.96100e-08 0.00000e+00 4.05500e-08 0.00000e+00
+ 4.05550e-08 2.00000e-03 4.06050e-08 2.00000e-03 4.06100e-08 0.00000e+00
+ 4.35500e-08 0.00000e+00 4.35550e-08 2.00000e-03 4.36050e-08 2.00000e-03
+ 4.36100e-08 0.00000e+00 4.45500e-08 0.00000e+00 4.45550e-08 2.00000e-03
+ 4.46050e-08 2.00000e-03 4.46100e-08 0.00000e+00 4.75500e-08 0.00000e+00
+ 4.75550e-08 2.00000e-03 4.76050e-08 2.00000e-03 4.76100e-08 0.00000e+00
+ 4.85500e-08 0.00000e+00 4.85550e-08 2.00000e-03 4.86050e-08 2.00000e-03
+ 4.86100e-08 0.00000e+00 5.15500e-08 0.00000e+00 5.15550e-08 2.00000e-03
+ 5.16050e-08 2.00000e-03 5.16100e-08 0.00000e+00 5.25500e-08 0.00000e+00
+ 5.25550e-08 2.00000e-03 5.26050e-08 2.00000e-03 5.26100e-08 0.00000e+00
+ 5.55500e-08 0.00000e+00 5.55550e-08 2.00000e-03 5.56050e-08 2.00000e-03
+ 5.56100e-08 0.00000e+00 5.65500e-08 0.00000e+00 5.65550e-08 2.00000e-03
+ 5.66050e-08 2.00000e-03 5.66100e-08 0.00000e+00 5.95500e-08 0.00000e+00
+ 5.95550e-08 2.00000e-03 5.96050e-08 2.00000e-03 5.96100e-08 0.00000e+00
+ 6.05500e-08 0.00000e+00 6.05550e-08 2.00000e-03 6.06050e-08 2.00000e-03
+ 6.06100e-08 0.00000e+00 6.35500e-08 0.00000e+00 6.35550e-08 2.00000e-03
+ 6.36050e-08 2.00000e-03 6.36100e-08 0.00000e+00 6.45500e-08 0.00000e+00
+ 6.45550e-08 2.00000e-03 6.46050e-08 2.00000e-03 6.46100e-08 0.00000e+00
+ 6.75500e-08 0.00000e+00 6.75550e-08 2.00000e-03 6.76050e-08 2.00000e-03
+ 6.76100e-08 0.00000e+00 6.85500e-08 0.00000e+00 6.85550e-08 2.00000e-03
+ 6.86050e-08 2.00000e-03 6.86100e-08 0.00000e+00 7.15500e-08 0.00000e+00
+ 7.15550e-08 2.00000e-03 7.16050e-08 2.00000e-03 7.16100e-08 0.00000e+00
+ 7.25500e-08 0.00000e+00 7.25550e-08 2.00000e-03 7.26050e-08 2.00000e-03
+ 7.26100e-08 0.00000e+00 7.55500e-08 0.00000e+00 7.55550e-08 2.00000e-03
+ 7.56050e-08 2.00000e-03 7.56100e-08 0.00000e+00 7.65500e-08 0.00000e+00
+ 7.65550e-08 2.00000e-03 7.66050e-08 2.00000e-03 7.66100e-08 0.00000e+00
+ 7.95500e-08 0.00000e+00 7.95550e-08 2.00000e-03 7.96050e-08 2.00000e-03
+ 7.96100e-08 0.00000e+00 8.05500e-08 0.00000e+00 8.05550e-08 2.00000e-03
+ 8.06050e-08 2.00000e-03 8.06100e-08 0.00000e+00 8.35500e-08 0.00000e+00
+ 8.35550e-08 2.00000e-03 8.36050e-08 2.00000e-03 8.36100e-08 0.00000e+00
+ 8.45500e-08 0.00000e+00 8.45550e-08 2.00000e-03 8.46050e-08 2.00000e-03
+ 8.46100e-08 0.00000e+00 8.75500e-08 0.00000e+00 8.75550e-08 2.00000e-03
+ 8.76050e-08 2.00000e-03 8.76100e-08 0.00000e+00 8.85500e-08 0.00000e+00
+ 8.85550e-08 2.00000e-03 8.86050e-08 2.00000e-03 8.86100e-08 0.00000e+00
+ 9.15500e-08 0.00000e+00 9.15550e-08 2.00000e-03 9.16050e-08 2.00000e-03
+ 9.16100e-08 0.00000e+00 9.25500e-08 0.00000e+00 9.25550e-08 2.00000e-03
+ 9.26050e-08 2.00000e-03 9.26100e-08 0.00000e+00 9.55500e-08 0.00000e+00
+ 9.55550e-08 2.00000e-03 9.56050e-08 2.00000e-03 9.56100e-08 0.00000e+00
+ 9.65500e-08 0.00000e+00 9.65550e-08 2.00000e-03 9.66050e-08 2.00000e-03
+ 9.66100e-08 0.00000e+00 9.95500e-08 0.00000e+00 9.95550e-08 2.00000e-03
+ 9.96050e-08 2.00000e-03 9.96100e-08 0.00000e+00 1.00550e-07 0.00000e+00
+ 1.00555e-07 2.00000e-03 1.00605e-07 2.00000e-03 1.00610e-07 0.00000e+00
+ 1.03550e-07 0.00000e+00 1.03555e-07 2.00000e-03 1.03605e-07 2.00000e-03
+ 1.03610e-07 0.00000e+00 1.04550e-07 0.00000e+00 1.04555e-07 2.00000e-03
+ 1.04605e-07 2.00000e-03 1.04610e-07 0.00000e+00 1.07550e-07 0.00000e+00
+ 1.07555e-07 2.00000e-03 1.07605e-07 2.00000e-03 1.07610e-07 0.00000e+00
+ 1.08550e-07 0.00000e+00 1.08555e-07 2.00000e-03 1.08605e-07 2.00000e-03
+ 1.08610e-07 0.00000e+00 1.11550e-07 0.00000e+00 1.11555e-07 2.00000e-03
+ 1.11605e-07 2.00000e-03 1.11610e-07 0.00000e+00 1.12550e-07 0.00000e+00
+ 1.12555e-07 2.00000e-03 1.12605e-07 2.00000e-03 1.12610e-07 0.00000e+00
+ 1.15550e-07 0.00000e+00 1.15555e-07 2.00000e-03 1.15605e-07 2.00000e-03
+ 1.15610e-07 0.00000e+00 1.16550e-07 0.00000e+00 1.16555e-07 2.00000e-03
+ 1.16605e-07 2.00000e-03 1.16610e-07 0.00000e+00 1.19550e-07 0.00000e+00
+ 1.19555e-07 2.00000e-03 1.19605e-07 2.00000e-03 1.19610e-07 0.00000e+00
+ 1.20550e-07 0.00000e+00 1.20555e-07 2.00000e-03 1.20605e-07 2.00000e-03
+ 1.20610e-07 0.00000e+00 1.23550e-07 0.00000e+00 1.23555e-07 2.00000e-03
+ 1.23605e-07 2.00000e-03 1.23610e-07 0.00000e+00 1.24550e-07 0.00000e+00
+ 1.24555e-07 2.00000e-03 1.24605e-07 2.00000e-03 1.24610e-07 0.00000e+00
+ 1.27550e-07 0.00000e+00 1.27555e-07 2.00000e-03 1.27605e-07 2.00000e-03
+ 1.27610e-07 0.00000e+00 1.28550e-07 0.00000e+00 1.28555e-07 2.00000e-03
+ 1.28605e-07 2.00000e-03 1.28610e-07 0.00000e+00 1.31550e-07 0.00000e+00
+ 1.31555e-07 2.00000e-03 1.31605e-07 2.00000e-03 1.31610e-07 0.00000e+00
+ 1.32550e-07 0.00000e+00 1.32555e-07 2.00000e-03 1.32605e-07 2.00000e-03
+ 1.32610e-07 0.00000e+00 1.35550e-07 0.00000e+00 1.35555e-07 2.00000e-03
+ 1.35605e-07 2.00000e-03 1.35610e-07 0.00000e+00 1.36550e-07 0.00000e+00
+ 1.36555e-07 2.00000e-03 1.36605e-07 2.00000e-03 1.36610e-07 0.00000e+00
+ 1.39550e-07 0.00000e+00 1.39555e-07 2.00000e-03 1.39605e-07 2.00000e-03
+ 1.39610e-07 0.00000e+00 1.40550e-07 0.00000e+00 1.40555e-07 2.00000e-03
+ 1.40605e-07 2.00000e-03 1.40610e-07 0.00000e+00 1.43550e-07 0.00000e+00
+ 1.43555e-07 2.00000e-03 1.43605e-07 2.00000e-03 1.43610e-07 0.00000e+00
+ 1.44550e-07 0.00000e+00 1.44555e-07 2.00000e-03 1.44605e-07 2.00000e-03
+ 1.44610e-07 0.00000e+00 1.47550e-07 0.00000e+00 1.47555e-07 2.00000e-03
+ 1.47605e-07 2.00000e-03 1.47610e-07 0.00000e+00 1.48550e-07 0.00000e+00
+ 1.48555e-07 2.00000e-03 1.48605e-07 2.00000e-03 1.48610e-07 0.00000e+00
+ 1.51550e-07 0.00000e+00 1.51555e-07 2.00000e-03 1.51605e-07 2.00000e-03
+ 1.51610e-07 0.00000e+00 1.52550e-07 0.00000e+00 1.52555e-07 2.00000e-03
+ 1.52605e-07 2.00000e-03 1.52610e-07 0.00000e+00 1.55550e-07 0.00000e+00
+ 1.55555e-07 2.00000e-03 1.55605e-07 2.00000e-03 1.55610e-07 0.00000e+00
+ 1.56550e-07 0.00000e+00 1.56555e-07 2.00000e-03 1.56605e-07 2.00000e-03
+ 1.56610e-07 0.00000e+00 1.59550e-07 0.00000e+00 1.59555e-07 2.00000e-03
+ 1.59605e-07 2.00000e-03 1.59610e-07 0.00000e+00 1.60550e-07 0.00000e+00
+ 1.60555e-07 2.00000e-03 1.60605e-07 2.00000e-03 1.60610e-07 0.00000e+00
+ 1.63550e-07 0.00000e+00 1.63555e-07 2.00000e-03 1.63605e-07 2.00000e-03
+ 1.63610e-07 0.00000e+00 1.64550e-07 0.00000e+00 1.64555e-07 2.00000e-03
+ 1.64605e-07 2.00000e-03 1.64610e-07 0.00000e+00 1.67550e-07 0.00000e+00
+ 1.67555e-07 2.00000e-03 1.67605e-07 2.00000e-03 1.67610e-07 0.00000e+00
+ 1.68550e-07 0.00000e+00 1.68555e-07 2.00000e-03 1.68605e-07 2.00000e-03
+ 1.68610e-07 0.00000e+00 1.71550e-07 0.00000e+00 1.71555e-07 2.00000e-03
+ 1.71605e-07 2.00000e-03 1.71610e-07 0.00000e+00 1.72550e-07 0.00000e+00
+ 1.72555e-07 2.00000e-03 1.72605e-07 2.00000e-03 1.72610e-07 0.00000e+00
+ 1.75550e-07 0.00000e+00 1.75555e-07 2.00000e-03 1.75605e-07 2.00000e-03
+ 1.75610e-07 0.00000e+00 1.76550e-07 0.00000e+00 1.76555e-07 2.00000e-03
+ 1.76605e-07 2.00000e-03 1.76610e-07 0.00000e+00 1.79550e-07 0.00000e+00
+ 1.79555e-07 2.00000e-03 1.79605e-07 2.00000e-03 1.79610e-07 0.00000e+00
+ 1.80550e-07 0.00000e+00 1.80555e-07 2.00000e-03 1.80605e-07 2.00000e-03
+ 1.80610e-07 0.00000e+00 1.83550e-07 0.00000e+00 1.83555e-07 2.00000e-03
+ 1.83605e-07 2.00000e-03 1.83610e-07 0.00000e+00 1.84550e-07 0.00000e+00
+ 1.84555e-07 2.00000e-03 1.84605e-07 2.00000e-03 1.84610e-07 0.00000e+00
+ 1.87550e-07 0.00000e+00 1.87555e-07 2.00000e-03 1.87605e-07 2.00000e-03
+ 1.87610e-07 0.00000e+00 1.88550e-07 0.00000e+00 1.88555e-07 2.00000e-03
+ 1.88605e-07 2.00000e-03 1.88610e-07 0.00000e+00 1.91550e-07 0.00000e+00
+ 1.91555e-07 2.00000e-03 1.91605e-07 2.00000e-03 1.91610e-07 0.00000e+00
+ 1.92550e-07 0.00000e+00 1.92555e-07 2.00000e-03 1.92605e-07 2.00000e-03
+ 1.92610e-07 0.00000e+00 1.95550e-07 0.00000e+00 1.95555e-07 2.00000e-03
+ 1.95605e-07 2.00000e-03 1.95610e-07 0.00000e+00 1.96550e-07 0.00000e+00
+ 1.96555e-07 2.00000e-03 1.96605e-07 2.00000e-03 1.96610e-07 0.00000e+00
+ 1.99550e-07 0.00000e+00 1.99555e-07 2.00000e-03 1.99605e-07 2.00000e-03
+ 1.99610e-07 0.00000e+00)
Iactualsynbias21 0 ACTUALSYNB21x PWL(0 0 7.40000e-10 0.00000e+00 7.65000e-10 6.70000e-04 8.00000e-10 0.00000e+00
+ 9.40000e-10 0.00000e+00 9.65000e-10 6.70000e-04 1.00000e-09 0.00000e+00
+ 1.14000e-09 0.00000e+00 1.16500e-09 6.70000e-04 1.20000e-09 0.00000e+00
+ 1.34000e-09 0.00000e+00 1.36500e-09 6.70000e-04 1.40000e-09 0.00000e+00
+ 1.54000e-09 0.00000e+00 1.56500e-09 6.70000e-04 1.60000e-09 0.00000e+00
+ 1.74000e-09 0.00000e+00 1.76500e-09 6.70000e-04 1.80000e-09 0.00000e+00
+ 1.94000e-09 0.00000e+00 1.96500e-09 6.70000e-04 2.00000e-09 0.00000e+00
+ 2.14000e-09 0.00000e+00 2.16500e-09 6.70000e-04 2.20000e-09 0.00000e+00
+ 2.34000e-09 0.00000e+00 2.36500e-09 6.70000e-04 2.40000e-09 0.00000e+00
+ 2.54000e-09 0.00000e+00 2.56500e-09 6.70000e-04 2.60000e-09 0.00000e+00
+ 2.74000e-09 0.00000e+00 2.76500e-09 6.70000e-04 2.80000e-09 0.00000e+00
+ 2.94000e-09 0.00000e+00 2.96500e-09 6.70000e-04 3.00000e-09 0.00000e+00
+ 3.14000e-09 0.00000e+00 3.16500e-09 6.70000e-04 3.20000e-09 0.00000e+00
+ 3.34000e-09 0.00000e+00 3.36500e-09 6.70000e-04 3.40000e-09 0.00000e+00
+ 3.54000e-09 0.00000e+00 3.56500e-09 6.70000e-04 3.60000e-09 0.00000e+00
+ 3.74000e-09 0.00000e+00 3.76500e-09 6.70000e-04 3.80000e-09 0.00000e+00
+ 3.94000e-09 0.00000e+00 3.96500e-09 6.70000e-04 4.00000e-09 0.00000e+00
+ 4.14000e-09 0.00000e+00 4.16500e-09 6.70000e-04 4.20000e-09 0.00000e+00
+ 4.34000e-09 0.00000e+00 4.36500e-09 6.70000e-04 4.40000e-09 0.00000e+00
+ 4.54000e-09 0.00000e+00 4.56500e-09 6.70000e-04 4.60000e-09 0.00000e+00
+ 4.74000e-09 0.00000e+00 4.76500e-09 6.70000e-04 4.80000e-09 0.00000e+00
+ 4.94000e-09 0.00000e+00 4.96500e-09 6.70000e-04 5.00000e-09 0.00000e+00
+ 5.14000e-09 0.00000e+00 5.16500e-09 6.70000e-04 5.20000e-09 0.00000e+00
+ 5.34000e-09 0.00000e+00 5.36500e-09 6.70000e-04 5.40000e-09 0.00000e+00
+ 5.54000e-09 0.00000e+00 5.56500e-09 6.70000e-04 5.60000e-09 0.00000e+00
+ 5.74000e-09 0.00000e+00 5.76500e-09 6.70000e-04 5.80000e-09 0.00000e+00
+ 5.94000e-09 0.00000e+00 5.96500e-09 6.70000e-04 6.00000e-09 0.00000e+00
+ 6.14000e-09 0.00000e+00 6.16500e-09 6.70000e-04 6.20000e-09 0.00000e+00
+ 6.34000e-09 0.00000e+00 6.36500e-09 6.70000e-04 6.40000e-09 0.00000e+00
+ 6.54000e-09 0.00000e+00 6.56500e-09 6.70000e-04 6.60000e-09 0.00000e+00
+ 6.74000e-09 0.00000e+00 6.76500e-09 6.70000e-04 6.80000e-09 0.00000e+00
+ 6.94000e-09 0.00000e+00 6.96500e-09 6.70000e-04 7.00000e-09 0.00000e+00
+ 7.14000e-09 0.00000e+00 7.16500e-09 6.70000e-04 7.20000e-09 0.00000e+00
+ 7.34000e-09 0.00000e+00 7.36500e-09 6.70000e-04 7.40000e-09 0.00000e+00
+ 7.54000e-09 0.00000e+00 7.56500e-09 6.70000e-04 7.60000e-09 0.00000e+00
+ 7.74000e-09 0.00000e+00 7.76500e-09 6.70000e-04 7.80000e-09 0.00000e+00
+ 7.94000e-09 0.00000e+00 7.96500e-09 6.70000e-04 8.00000e-09 0.00000e+00
+ 8.14000e-09 0.00000e+00 8.16500e-09 6.70000e-04 8.20000e-09 0.00000e+00
+ 8.34000e-09 0.00000e+00 8.36500e-09 6.70000e-04 8.40000e-09 0.00000e+00
+ 8.54000e-09 0.00000e+00 8.56500e-09 6.70000e-04 8.60000e-09 0.00000e+00
+ 8.74000e-09 0.00000e+00 8.76500e-09 6.70000e-04 8.80000e-09 0.00000e+00
+ 8.94000e-09 0.00000e+00 8.96500e-09 6.70000e-04 9.00000e-09 0.00000e+00
+ 9.14000e-09 0.00000e+00 9.16500e-09 6.70000e-04 9.20000e-09 0.00000e+00
+ 9.34000e-09 0.00000e+00 9.36500e-09 6.70000e-04 9.40000e-09 0.00000e+00
+ 9.54000e-09 0.00000e+00 9.56500e-09 6.70000e-04 9.60000e-09 0.00000e+00
+ 9.74000e-09 0.00000e+00 9.76500e-09 6.70000e-04 9.80000e-09 0.00000e+00
+ 9.94000e-09 0.00000e+00 9.96500e-09 6.70000e-04 1.00000e-08 0.00000e+00
+ 1.01400e-08 0.00000e+00 1.01650e-08 6.70000e-04 1.02000e-08 0.00000e+00
+ 1.03400e-08 0.00000e+00 1.03650e-08 6.70000e-04 1.04000e-08 0.00000e+00
+ 1.05400e-08 0.00000e+00 1.05650e-08 6.70000e-04 1.06000e-08 0.00000e+00
+ 1.07400e-08 0.00000e+00 1.07650e-08 6.70000e-04 1.08000e-08 0.00000e+00
+ 1.09400e-08 0.00000e+00 1.09650e-08 6.70000e-04 1.10000e-08 0.00000e+00
+ 1.11400e-08 0.00000e+00 1.11650e-08 6.70000e-04 1.12000e-08 0.00000e+00
+ 1.13400e-08 0.00000e+00 1.13650e-08 6.70000e-04 1.14000e-08 0.00000e+00
+ 1.15400e-08 0.00000e+00 1.15650e-08 6.70000e-04 1.16000e-08 0.00000e+00
+ 1.17400e-08 0.00000e+00 1.17650e-08 6.70000e-04 1.18000e-08 0.00000e+00
+ 1.19400e-08 0.00000e+00 1.19650e-08 6.70000e-04 1.20000e-08 0.00000e+00
+ 1.21400e-08 0.00000e+00 1.21650e-08 6.70000e-04 1.22000e-08 0.00000e+00
+ 1.23400e-08 0.00000e+00 1.23650e-08 6.70000e-04 1.24000e-08 0.00000e+00
+ 1.25400e-08 0.00000e+00 1.25650e-08 6.70000e-04 1.26000e-08 0.00000e+00
+ 1.27400e-08 0.00000e+00 1.27650e-08 6.70000e-04 1.28000e-08 0.00000e+00
+ 1.29400e-08 0.00000e+00 1.29650e-08 6.70000e-04 1.30000e-08 0.00000e+00
+ 1.31400e-08 0.00000e+00 1.31650e-08 6.70000e-04 1.32000e-08 0.00000e+00
+ 1.33400e-08 0.00000e+00 1.33650e-08 6.70000e-04 1.34000e-08 0.00000e+00
+ 1.35400e-08 0.00000e+00 1.35650e-08 6.70000e-04 1.36000e-08 0.00000e+00
+ 1.37400e-08 0.00000e+00 1.37650e-08 6.70000e-04 1.38000e-08 0.00000e+00
+ 1.39400e-08 0.00000e+00 1.39650e-08 6.70000e-04 1.40000e-08 0.00000e+00
+ 1.41400e-08 0.00000e+00 1.41650e-08 6.70000e-04 1.42000e-08 0.00000e+00
+ 1.43400e-08 0.00000e+00 1.43650e-08 6.70000e-04 1.44000e-08 0.00000e+00
+ 1.45400e-08 0.00000e+00 1.45650e-08 6.70000e-04 1.46000e-08 0.00000e+00
+ 1.47400e-08 0.00000e+00 1.47650e-08 6.70000e-04 1.48000e-08 0.00000e+00
+ 1.49400e-08 0.00000e+00 1.49650e-08 6.70000e-04 1.50000e-08 0.00000e+00
+ 1.51400e-08 0.00000e+00 1.51650e-08 6.70000e-04 1.52000e-08 0.00000e+00
+ 1.53400e-08 0.00000e+00 1.53650e-08 6.70000e-04 1.54000e-08 0.00000e+00
+ 1.55400e-08 0.00000e+00 1.55650e-08 6.70000e-04 1.56000e-08 0.00000e+00
+ 1.57400e-08 0.00000e+00 1.57650e-08 6.70000e-04 1.58000e-08 0.00000e+00
+ 1.59400e-08 0.00000e+00 1.59650e-08 6.70000e-04 1.60000e-08 0.00000e+00
+ 1.61400e-08 0.00000e+00 1.61650e-08 6.70000e-04 1.62000e-08 0.00000e+00
+ 1.63400e-08 0.00000e+00 1.63650e-08 6.70000e-04 1.64000e-08 0.00000e+00
+ 1.65400e-08 0.00000e+00 1.65650e-08 6.70000e-04 1.66000e-08 0.00000e+00
+ 1.67400e-08 0.00000e+00 1.67650e-08 6.70000e-04 1.68000e-08 0.00000e+00
+ 1.69400e-08 0.00000e+00 1.69650e-08 6.70000e-04 1.70000e-08 0.00000e+00
+ 1.71400e-08 0.00000e+00 1.71650e-08 6.70000e-04 1.72000e-08 0.00000e+00
+ 1.73400e-08 0.00000e+00 1.73650e-08 6.70000e-04 1.74000e-08 0.00000e+00
+ 1.75400e-08 0.00000e+00 1.75650e-08 6.70000e-04 1.76000e-08 0.00000e+00
+ 1.77400e-08 0.00000e+00 1.77650e-08 6.70000e-04 1.78000e-08 0.00000e+00
+ 1.79400e-08 0.00000e+00 1.79650e-08 6.70000e-04 1.80000e-08 0.00000e+00
+ 1.81400e-08 0.00000e+00 1.81650e-08 6.70000e-04 1.82000e-08 0.00000e+00
+ 1.83400e-08 0.00000e+00 1.83650e-08 6.70000e-04 1.84000e-08 0.00000e+00
+ 1.85400e-08 0.00000e+00 1.85650e-08 6.70000e-04 1.86000e-08 0.00000e+00
+ 1.87400e-08 0.00000e+00 1.87650e-08 6.70000e-04 1.88000e-08 0.00000e+00
+ 1.89400e-08 0.00000e+00 1.89650e-08 6.70000e-04 1.90000e-08 0.00000e+00
+ 1.91400e-08 0.00000e+00 1.91650e-08 6.70000e-04 1.92000e-08 0.00000e+00
+ 1.93400e-08 0.00000e+00 1.93650e-08 6.70000e-04 1.94000e-08 0.00000e+00
+ 1.95400e-08 0.00000e+00 1.95650e-08 6.70000e-04 1.96000e-08 0.00000e+00
+ 1.97400e-08 0.00000e+00 1.97650e-08 6.70000e-04 1.98000e-08 0.00000e+00
+ 1.99400e-08 0.00000e+00 1.99650e-08 6.70000e-04 2.00000e-08 0.00000e+00
+ 2.01400e-08 0.00000e+00 2.01650e-08 6.70000e-04 2.02000e-08 0.00000e+00
+ 2.03400e-08 0.00000e+00 2.03650e-08 6.70000e-04 2.04000e-08 0.00000e+00
+ 2.05400e-08 0.00000e+00 2.05650e-08 6.70000e-04 2.06000e-08 0.00000e+00
+ 2.07400e-08 0.00000e+00 2.07650e-08 6.70000e-04 2.08000e-08 0.00000e+00
+ 2.09400e-08 0.00000e+00 2.09650e-08 6.70000e-04 2.10000e-08 0.00000e+00
+ 2.11400e-08 0.00000e+00 2.11650e-08 6.70000e-04 2.12000e-08 0.00000e+00
+ 2.13400e-08 0.00000e+00 2.13650e-08 6.70000e-04 2.14000e-08 0.00000e+00
+ 2.15400e-08 0.00000e+00 2.15650e-08 6.70000e-04 2.16000e-08 0.00000e+00
+ 2.17400e-08 0.00000e+00 2.17650e-08 6.70000e-04 2.18000e-08 0.00000e+00
+ 2.19400e-08 0.00000e+00 2.19650e-08 6.70000e-04 2.20000e-08 0.00000e+00
+ 2.21400e-08 0.00000e+00 2.21650e-08 6.70000e-04 2.22000e-08 0.00000e+00
+ 2.23400e-08 0.00000e+00 2.23650e-08 6.70000e-04 2.24000e-08 0.00000e+00
+ 2.25400e-08 0.00000e+00 2.25650e-08 6.70000e-04 2.26000e-08 0.00000e+00
+ 2.27400e-08 0.00000e+00 2.27650e-08 6.70000e-04 2.28000e-08 0.00000e+00
+ 2.29400e-08 0.00000e+00 2.29650e-08 6.70000e-04 2.30000e-08 0.00000e+00
+ 2.31400e-08 0.00000e+00 2.31650e-08 6.70000e-04 2.32000e-08 0.00000e+00
+ 2.33400e-08 0.00000e+00 2.33650e-08 6.70000e-04 2.34000e-08 0.00000e+00
+ 2.35400e-08 0.00000e+00 2.35650e-08 6.70000e-04 2.36000e-08 0.00000e+00
+ 2.37400e-08 0.00000e+00 2.37650e-08 6.70000e-04 2.38000e-08 0.00000e+00
+ 2.39400e-08 0.00000e+00 2.39650e-08 6.70000e-04 2.40000e-08 0.00000e+00
+ 2.41400e-08 0.00000e+00 2.41650e-08 6.70000e-04 2.42000e-08 0.00000e+00
+ 2.43400e-08 0.00000e+00 2.43650e-08 6.70000e-04 2.44000e-08 0.00000e+00
+ 2.45400e-08 0.00000e+00 2.45650e-08 6.70000e-04 2.46000e-08 0.00000e+00
+ 2.47400e-08 0.00000e+00 2.47650e-08 6.70000e-04 2.48000e-08 0.00000e+00
+ 2.49400e-08 0.00000e+00 2.49650e-08 6.70000e-04 2.50000e-08 0.00000e+00
+ 2.51400e-08 0.00000e+00 2.51650e-08 6.70000e-04 2.52000e-08 0.00000e+00
+ 2.53400e-08 0.00000e+00 2.53650e-08 6.70000e-04 2.54000e-08 0.00000e+00
+ 2.55400e-08 0.00000e+00 2.55650e-08 6.70000e-04 2.56000e-08 0.00000e+00
+ 2.57400e-08 0.00000e+00 2.57650e-08 6.70000e-04 2.58000e-08 0.00000e+00
+ 2.59400e-08 0.00000e+00 2.59650e-08 6.70000e-04 2.60000e-08 0.00000e+00
+ 2.61400e-08 0.00000e+00 2.61650e-08 6.70000e-04 2.62000e-08 0.00000e+00
+ 2.63400e-08 0.00000e+00 2.63650e-08 6.70000e-04 2.64000e-08 0.00000e+00
+ 2.65400e-08 0.00000e+00 2.65650e-08 6.70000e-04 2.66000e-08 0.00000e+00
+ 2.67400e-08 0.00000e+00 2.67650e-08 6.70000e-04 2.68000e-08 0.00000e+00
+ 2.69400e-08 0.00000e+00 2.69650e-08 6.70000e-04 2.70000e-08 0.00000e+00
+ 2.71400e-08 0.00000e+00 2.71650e-08 6.70000e-04 2.72000e-08 0.00000e+00
+ 2.73400e-08 0.00000e+00 2.73650e-08 6.70000e-04 2.74000e-08 0.00000e+00
+ 2.75400e-08 0.00000e+00 2.75650e-08 6.70000e-04 2.76000e-08 0.00000e+00
+ 2.77400e-08 0.00000e+00 2.77650e-08 6.70000e-04 2.78000e-08 0.00000e+00
+ 2.79400e-08 0.00000e+00 2.79650e-08 6.70000e-04 2.80000e-08 0.00000e+00
+ 2.81400e-08 0.00000e+00 2.81650e-08 6.70000e-04 2.82000e-08 0.00000e+00
+ 2.83400e-08 0.00000e+00 2.83650e-08 6.70000e-04 2.84000e-08 0.00000e+00
+ 2.85400e-08 0.00000e+00 2.85650e-08 6.70000e-04 2.86000e-08 0.00000e+00
+ 2.87400e-08 0.00000e+00 2.87650e-08 6.70000e-04 2.88000e-08 0.00000e+00
+ 2.89400e-08 0.00000e+00 2.89650e-08 6.70000e-04 2.90000e-08 0.00000e+00
+ 2.91400e-08 0.00000e+00 2.91650e-08 6.70000e-04 2.92000e-08 0.00000e+00
+ 2.93400e-08 0.00000e+00 2.93650e-08 6.70000e-04 2.94000e-08 0.00000e+00
+ 2.95400e-08 0.00000e+00 2.95650e-08 6.70000e-04 2.96000e-08 0.00000e+00
+ 2.97400e-08 0.00000e+00 2.97650e-08 6.70000e-04 2.98000e-08 0.00000e+00
+ 2.99400e-08 0.00000e+00 2.99650e-08 6.70000e-04 3.00000e-08 0.00000e+00
+ 3.01400e-08 0.00000e+00 3.01650e-08 6.70000e-04 3.02000e-08 0.00000e+00
+ 3.03400e-08 0.00000e+00 3.03650e-08 6.70000e-04 3.04000e-08 0.00000e+00
+ 3.05400e-08 0.00000e+00 3.05650e-08 6.70000e-04 3.06000e-08 0.00000e+00
+ 3.07400e-08 0.00000e+00 3.07650e-08 6.70000e-04 3.08000e-08 0.00000e+00
+ 3.09400e-08 0.00000e+00 3.09650e-08 6.70000e-04 3.10000e-08 0.00000e+00
+ 3.11400e-08 0.00000e+00 3.11650e-08 6.70000e-04 3.12000e-08 0.00000e+00
+ 3.13400e-08 0.00000e+00 3.13650e-08 6.70000e-04 3.14000e-08 0.00000e+00
+ 3.15400e-08 0.00000e+00 3.15650e-08 6.70000e-04 3.16000e-08 0.00000e+00
+ 3.17400e-08 0.00000e+00 3.17650e-08 6.70000e-04 3.18000e-08 0.00000e+00
+ 3.19400e-08 0.00000e+00 3.19650e-08 6.70000e-04 3.20000e-08 0.00000e+00
+ 3.21400e-08 0.00000e+00 3.21650e-08 6.70000e-04 3.22000e-08 0.00000e+00
+ 3.23400e-08 0.00000e+00 3.23650e-08 6.70000e-04 3.24000e-08 0.00000e+00
+ 3.25400e-08 0.00000e+00 3.25650e-08 6.70000e-04 3.26000e-08 0.00000e+00
+ 3.27400e-08 0.00000e+00 3.27650e-08 6.70000e-04 3.28000e-08 0.00000e+00
+ 3.29400e-08 0.00000e+00 3.29650e-08 6.70000e-04 3.30000e-08 0.00000e+00
+ 3.31400e-08 0.00000e+00 3.31650e-08 6.70000e-04 3.32000e-08 0.00000e+00
+ 3.33400e-08 0.00000e+00 3.33650e-08 6.70000e-04 3.34000e-08 0.00000e+00
+ 3.35400e-08 0.00000e+00 3.35650e-08 6.70000e-04 3.36000e-08 0.00000e+00
+ 3.37400e-08 0.00000e+00 3.37650e-08 6.70000e-04 3.38000e-08 0.00000e+00
+ 3.39400e-08 0.00000e+00 3.39650e-08 6.70000e-04 3.40000e-08 0.00000e+00
+ 3.41400e-08 0.00000e+00 3.41650e-08 6.70000e-04 3.42000e-08 0.00000e+00
+ 3.43400e-08 0.00000e+00 3.43650e-08 6.70000e-04 3.44000e-08 0.00000e+00
+ 3.45400e-08 0.00000e+00 3.45650e-08 6.70000e-04 3.46000e-08 0.00000e+00
+ 3.47400e-08 0.00000e+00 3.47650e-08 6.70000e-04 3.48000e-08 0.00000e+00
+ 3.49400e-08 0.00000e+00 3.49650e-08 6.70000e-04 3.50000e-08 0.00000e+00
+ 3.51400e-08 0.00000e+00 3.51650e-08 6.70000e-04 3.52000e-08 0.00000e+00
+ 3.53400e-08 0.00000e+00 3.53650e-08 6.70000e-04 3.54000e-08 0.00000e+00
+ 3.55400e-08 0.00000e+00 3.55650e-08 6.70000e-04 3.56000e-08 0.00000e+00
+ 3.57400e-08 0.00000e+00 3.57650e-08 6.70000e-04 3.58000e-08 0.00000e+00
+ 3.59400e-08 0.00000e+00 3.59650e-08 6.70000e-04 3.60000e-08 0.00000e+00
+ 3.61400e-08 0.00000e+00 3.61650e-08 6.70000e-04 3.62000e-08 0.00000e+00
+ 3.63400e-08 0.00000e+00 3.63650e-08 6.70000e-04 3.64000e-08 0.00000e+00
+ 3.65400e-08 0.00000e+00 3.65650e-08 6.70000e-04 3.66000e-08 0.00000e+00
+ 3.67400e-08 0.00000e+00 3.67650e-08 6.70000e-04 3.68000e-08 0.00000e+00
+ 3.69400e-08 0.00000e+00 3.69650e-08 6.70000e-04 3.70000e-08 0.00000e+00
+ 3.71400e-08 0.00000e+00 3.71650e-08 6.70000e-04 3.72000e-08 0.00000e+00
+ 3.73400e-08 0.00000e+00 3.73650e-08 6.70000e-04 3.74000e-08 0.00000e+00
+ 3.75400e-08 0.00000e+00 3.75650e-08 6.70000e-04 3.76000e-08 0.00000e+00
+ 3.77400e-08 0.00000e+00 3.77650e-08 6.70000e-04 3.78000e-08 0.00000e+00
+ 3.79400e-08 0.00000e+00 3.79650e-08 6.70000e-04 3.80000e-08 0.00000e+00
+ 3.81400e-08 0.00000e+00 3.81650e-08 6.70000e-04 3.82000e-08 0.00000e+00
+ 3.83400e-08 0.00000e+00 3.83650e-08 6.70000e-04 3.84000e-08 0.00000e+00
+ 3.85400e-08 0.00000e+00 3.85650e-08 6.70000e-04 3.86000e-08 0.00000e+00
+ 3.87400e-08 0.00000e+00 3.87650e-08 6.70000e-04 3.88000e-08 0.00000e+00
+ 3.89400e-08 0.00000e+00 3.89650e-08 6.70000e-04 3.90000e-08 0.00000e+00
+ 3.91400e-08 0.00000e+00 3.91650e-08 6.70000e-04 3.92000e-08 0.00000e+00
+ 3.93400e-08 0.00000e+00 3.93650e-08 6.70000e-04 3.94000e-08 0.00000e+00
+ 3.95400e-08 0.00000e+00 3.95650e-08 6.70000e-04 3.96000e-08 0.00000e+00
+ 3.97400e-08 0.00000e+00 3.97650e-08 6.70000e-04 3.98000e-08 0.00000e+00
+ 3.99400e-08 0.00000e+00 3.99650e-08 6.70000e-04 4.00000e-08 0.00000e+00
+ 4.01400e-08 0.00000e+00 4.01650e-08 6.70000e-04 4.02000e-08 0.00000e+00
+ 4.03400e-08 0.00000e+00 4.03650e-08 6.70000e-04 4.04000e-08 0.00000e+00
+ 4.05400e-08 0.00000e+00 4.05650e-08 6.70000e-04 4.06000e-08 0.00000e+00
+ 4.07400e-08 0.00000e+00 4.07650e-08 6.70000e-04 4.08000e-08 0.00000e+00
+ 4.09400e-08 0.00000e+00 4.09650e-08 6.70000e-04 4.10000e-08 0.00000e+00
+ 4.11400e-08 0.00000e+00 4.11650e-08 6.70000e-04 4.12000e-08 0.00000e+00
+ 4.13400e-08 0.00000e+00 4.13650e-08 6.70000e-04 4.14000e-08 0.00000e+00
+ 4.15400e-08 0.00000e+00 4.15650e-08 6.70000e-04 4.16000e-08 0.00000e+00
+ 4.17400e-08 0.00000e+00 4.17650e-08 6.70000e-04 4.18000e-08 0.00000e+00
+ 4.19400e-08 0.00000e+00 4.19650e-08 6.70000e-04 4.20000e-08 0.00000e+00
+ 4.21400e-08 0.00000e+00 4.21650e-08 6.70000e-04 4.22000e-08 0.00000e+00
+ 4.23400e-08 0.00000e+00 4.23650e-08 6.70000e-04 4.24000e-08 0.00000e+00
+ 4.25400e-08 0.00000e+00 4.25650e-08 6.70000e-04 4.26000e-08 0.00000e+00
+ 4.27400e-08 0.00000e+00 4.27650e-08 6.70000e-04 4.28000e-08 0.00000e+00
+ 4.29400e-08 0.00000e+00 4.29650e-08 6.70000e-04 4.30000e-08 0.00000e+00
+ 4.31400e-08 0.00000e+00 4.31650e-08 6.70000e-04 4.32000e-08 0.00000e+00
+ 4.33400e-08 0.00000e+00 4.33650e-08 6.70000e-04 4.34000e-08 0.00000e+00
+ 4.35400e-08 0.00000e+00 4.35650e-08 6.70000e-04 4.36000e-08 0.00000e+00
+ 4.37400e-08 0.00000e+00 4.37650e-08 6.70000e-04 4.38000e-08 0.00000e+00
+ 4.39400e-08 0.00000e+00 4.39650e-08 6.70000e-04 4.40000e-08 0.00000e+00
+ 4.41400e-08 0.00000e+00 4.41650e-08 6.70000e-04 4.42000e-08 0.00000e+00
+ 4.43400e-08 0.00000e+00 4.43650e-08 6.70000e-04 4.44000e-08 0.00000e+00
+ 4.45400e-08 0.00000e+00 4.45650e-08 6.70000e-04 4.46000e-08 0.00000e+00
+ 4.47400e-08 0.00000e+00 4.47650e-08 6.70000e-04 4.48000e-08 0.00000e+00
+ 4.49400e-08 0.00000e+00 4.49650e-08 6.70000e-04 4.50000e-08 0.00000e+00
+ 4.51400e-08 0.00000e+00 4.51650e-08 6.70000e-04 4.52000e-08 0.00000e+00
+ 4.53400e-08 0.00000e+00 4.53650e-08 6.70000e-04 4.54000e-08 0.00000e+00
+ 4.55400e-08 0.00000e+00 4.55650e-08 6.70000e-04 4.56000e-08 0.00000e+00
+ 4.57400e-08 0.00000e+00 4.57650e-08 6.70000e-04 4.58000e-08 0.00000e+00
+ 4.59400e-08 0.00000e+00 4.59650e-08 6.70000e-04 4.60000e-08 0.00000e+00
+ 4.61400e-08 0.00000e+00 4.61650e-08 6.70000e-04 4.62000e-08 0.00000e+00
+ 4.63400e-08 0.00000e+00 4.63650e-08 6.70000e-04 4.64000e-08 0.00000e+00
+ 4.65400e-08 0.00000e+00 4.65650e-08 6.70000e-04 4.66000e-08 0.00000e+00
+ 4.67400e-08 0.00000e+00 4.67650e-08 6.70000e-04 4.68000e-08 0.00000e+00
+ 4.69400e-08 0.00000e+00 4.69650e-08 6.70000e-04 4.70000e-08 0.00000e+00
+ 4.71400e-08 0.00000e+00 4.71650e-08 6.70000e-04 4.72000e-08 0.00000e+00
+ 4.73400e-08 0.00000e+00 4.73650e-08 6.70000e-04 4.74000e-08 0.00000e+00
+ 4.75400e-08 0.00000e+00 4.75650e-08 6.70000e-04 4.76000e-08 0.00000e+00
+ 4.77400e-08 0.00000e+00 4.77650e-08 6.70000e-04 4.78000e-08 0.00000e+00
+ 4.79400e-08 0.00000e+00 4.79650e-08 6.70000e-04 4.80000e-08 0.00000e+00
+ 4.81400e-08 0.00000e+00 4.81650e-08 6.70000e-04 4.82000e-08 0.00000e+00
+ 4.83400e-08 0.00000e+00 4.83650e-08 6.70000e-04 4.84000e-08 0.00000e+00
+ 4.85400e-08 0.00000e+00 4.85650e-08 6.70000e-04 4.86000e-08 0.00000e+00
+ 4.87400e-08 0.00000e+00 4.87650e-08 6.70000e-04 4.88000e-08 0.00000e+00
+ 4.89400e-08 0.00000e+00 4.89650e-08 6.70000e-04 4.90000e-08 0.00000e+00
+ 4.91400e-08 0.00000e+00 4.91650e-08 6.70000e-04 4.92000e-08 0.00000e+00
+ 4.93400e-08 0.00000e+00 4.93650e-08 6.70000e-04 4.94000e-08 0.00000e+00
+ 4.95400e-08 0.00000e+00 4.95650e-08 6.70000e-04 4.96000e-08 0.00000e+00
+ 4.97400e-08 0.00000e+00 4.97650e-08 6.70000e-04 4.98000e-08 0.00000e+00
+ 4.99400e-08 0.00000e+00 4.99650e-08 6.70000e-04 5.00000e-08 0.00000e+00
+ 5.01400e-08 0.00000e+00 5.01650e-08 6.70000e-04 5.02000e-08 0.00000e+00
+ 5.03400e-08 0.00000e+00 5.03650e-08 6.70000e-04 5.04000e-08 0.00000e+00
+ 5.05400e-08 0.00000e+00 5.05650e-08 6.70000e-04 5.06000e-08 0.00000e+00
+ 5.07400e-08 0.00000e+00 5.07650e-08 6.70000e-04 5.08000e-08 0.00000e+00
+ 5.09400e-08 0.00000e+00 5.09650e-08 6.70000e-04 5.10000e-08 0.00000e+00
+ 5.11400e-08 0.00000e+00 5.11650e-08 6.70000e-04 5.12000e-08 0.00000e+00
+ 5.13400e-08 0.00000e+00 5.13650e-08 6.70000e-04 5.14000e-08 0.00000e+00
+ 5.15400e-08 0.00000e+00 5.15650e-08 6.70000e-04 5.16000e-08 0.00000e+00
+ 5.17400e-08 0.00000e+00 5.17650e-08 6.70000e-04 5.18000e-08 0.00000e+00
+ 5.19400e-08 0.00000e+00 5.19650e-08 6.70000e-04 5.20000e-08 0.00000e+00
+ 5.21400e-08 0.00000e+00 5.21650e-08 6.70000e-04 5.22000e-08 0.00000e+00
+ 5.23400e-08 0.00000e+00 5.23650e-08 6.70000e-04 5.24000e-08 0.00000e+00
+ 5.25400e-08 0.00000e+00 5.25650e-08 6.70000e-04 5.26000e-08 0.00000e+00
+ 5.27400e-08 0.00000e+00 5.27650e-08 6.70000e-04 5.28000e-08 0.00000e+00
+ 5.29400e-08 0.00000e+00 5.29650e-08 6.70000e-04 5.30000e-08 0.00000e+00
+ 5.31400e-08 0.00000e+00 5.31650e-08 6.70000e-04 5.32000e-08 0.00000e+00
+ 5.33400e-08 0.00000e+00 5.33650e-08 6.70000e-04 5.34000e-08 0.00000e+00
+ 5.35400e-08 0.00000e+00 5.35650e-08 6.70000e-04 5.36000e-08 0.00000e+00
+ 5.37400e-08 0.00000e+00 5.37650e-08 6.70000e-04 5.38000e-08 0.00000e+00
+ 5.39400e-08 0.00000e+00 5.39650e-08 6.70000e-04 5.40000e-08 0.00000e+00
+ 5.41400e-08 0.00000e+00 5.41650e-08 6.70000e-04 5.42000e-08 0.00000e+00
+ 5.43400e-08 0.00000e+00 5.43650e-08 6.70000e-04 5.44000e-08 0.00000e+00
+ 5.45400e-08 0.00000e+00 5.45650e-08 6.70000e-04 5.46000e-08 0.00000e+00
+ 5.47400e-08 0.00000e+00 5.47650e-08 6.70000e-04 5.48000e-08 0.00000e+00
+ 5.49400e-08 0.00000e+00 5.49650e-08 6.70000e-04 5.50000e-08 0.00000e+00
+ 5.51400e-08 0.00000e+00 5.51650e-08 6.70000e-04 5.52000e-08 0.00000e+00
+ 5.53400e-08 0.00000e+00 5.53650e-08 6.70000e-04 5.54000e-08 0.00000e+00
+ 5.55400e-08 0.00000e+00 5.55650e-08 6.70000e-04 5.56000e-08 0.00000e+00
+ 5.57400e-08 0.00000e+00 5.57650e-08 6.70000e-04 5.58000e-08 0.00000e+00
+ 5.59400e-08 0.00000e+00 5.59650e-08 6.70000e-04 5.60000e-08 0.00000e+00
+ 5.61400e-08 0.00000e+00 5.61650e-08 6.70000e-04 5.62000e-08 0.00000e+00
+ 5.63400e-08 0.00000e+00 5.63650e-08 6.70000e-04 5.64000e-08 0.00000e+00
+ 5.65400e-08 0.00000e+00 5.65650e-08 6.70000e-04 5.66000e-08 0.00000e+00
+ 5.67400e-08 0.00000e+00 5.67650e-08 6.70000e-04 5.68000e-08 0.00000e+00
+ 5.69400e-08 0.00000e+00 5.69650e-08 6.70000e-04 5.70000e-08 0.00000e+00
+ 5.71400e-08 0.00000e+00 5.71650e-08 6.70000e-04 5.72000e-08 0.00000e+00
+ 5.73400e-08 0.00000e+00 5.73650e-08 6.70000e-04 5.74000e-08 0.00000e+00
+ 5.75400e-08 0.00000e+00 5.75650e-08 6.70000e-04 5.76000e-08 0.00000e+00
+ 5.77400e-08 0.00000e+00 5.77650e-08 6.70000e-04 5.78000e-08 0.00000e+00
+ 5.79400e-08 0.00000e+00 5.79650e-08 6.70000e-04 5.80000e-08 0.00000e+00
+ 5.81400e-08 0.00000e+00 5.81650e-08 6.70000e-04 5.82000e-08 0.00000e+00
+ 5.83400e-08 0.00000e+00 5.83650e-08 6.70000e-04 5.84000e-08 0.00000e+00
+ 5.85400e-08 0.00000e+00 5.85650e-08 6.70000e-04 5.86000e-08 0.00000e+00
+ 5.87400e-08 0.00000e+00 5.87650e-08 6.70000e-04 5.88000e-08 0.00000e+00
+ 5.89400e-08 0.00000e+00 5.89650e-08 6.70000e-04 5.90000e-08 0.00000e+00
+ 5.91400e-08 0.00000e+00 5.91650e-08 6.70000e-04 5.92000e-08 0.00000e+00
+ 5.93400e-08 0.00000e+00 5.93650e-08 6.70000e-04 5.94000e-08 0.00000e+00
+ 5.95400e-08 0.00000e+00 5.95650e-08 6.70000e-04 5.96000e-08 0.00000e+00
+ 5.97400e-08 0.00000e+00 5.97650e-08 6.70000e-04 5.98000e-08 0.00000e+00
+ 5.99400e-08 0.00000e+00 5.99650e-08 6.70000e-04 6.00000e-08 0.00000e+00
+ 6.01400e-08 0.00000e+00 6.01650e-08 6.70000e-04 6.02000e-08 0.00000e+00
+ 6.03400e-08 0.00000e+00 6.03650e-08 6.70000e-04 6.04000e-08 0.00000e+00
+ 6.05400e-08 0.00000e+00 6.05650e-08 6.70000e-04 6.06000e-08 0.00000e+00
+ 6.07400e-08 0.00000e+00 6.07650e-08 6.70000e-04 6.08000e-08 0.00000e+00
+ 6.09400e-08 0.00000e+00 6.09650e-08 6.70000e-04 6.10000e-08 0.00000e+00
+ 6.11400e-08 0.00000e+00 6.11650e-08 6.70000e-04 6.12000e-08 0.00000e+00
+ 6.13400e-08 0.00000e+00 6.13650e-08 6.70000e-04 6.14000e-08 0.00000e+00
+ 6.15400e-08 0.00000e+00 6.15650e-08 6.70000e-04 6.16000e-08 0.00000e+00
+ 6.17400e-08 0.00000e+00 6.17650e-08 6.70000e-04 6.18000e-08 0.00000e+00
+ 6.19400e-08 0.00000e+00 6.19650e-08 6.70000e-04 6.20000e-08 0.00000e+00
+ 6.21400e-08 0.00000e+00 6.21650e-08 6.70000e-04 6.22000e-08 0.00000e+00
+ 6.23400e-08 0.00000e+00 6.23650e-08 6.70000e-04 6.24000e-08 0.00000e+00
+ 6.25400e-08 0.00000e+00 6.25650e-08 6.70000e-04 6.26000e-08 0.00000e+00
+ 6.27400e-08 0.00000e+00 6.27650e-08 6.70000e-04 6.28000e-08 0.00000e+00
+ 6.29400e-08 0.00000e+00 6.29650e-08 6.70000e-04 6.30000e-08 0.00000e+00
+ 6.31400e-08 0.00000e+00 6.31650e-08 6.70000e-04 6.32000e-08 0.00000e+00
+ 6.33400e-08 0.00000e+00 6.33650e-08 6.70000e-04 6.34000e-08 0.00000e+00
+ 6.35400e-08 0.00000e+00 6.35650e-08 6.70000e-04 6.36000e-08 0.00000e+00
+ 6.37400e-08 0.00000e+00 6.37650e-08 6.70000e-04 6.38000e-08 0.00000e+00
+ 6.39400e-08 0.00000e+00 6.39650e-08 6.70000e-04 6.40000e-08 0.00000e+00
+ 6.41400e-08 0.00000e+00 6.41650e-08 6.70000e-04 6.42000e-08 0.00000e+00
+ 6.43400e-08 0.00000e+00 6.43650e-08 6.70000e-04 6.44000e-08 0.00000e+00
+ 6.45400e-08 0.00000e+00 6.45650e-08 6.70000e-04 6.46000e-08 0.00000e+00
+ 6.47400e-08 0.00000e+00 6.47650e-08 6.70000e-04 6.48000e-08 0.00000e+00
+ 6.49400e-08 0.00000e+00 6.49650e-08 6.70000e-04 6.50000e-08 0.00000e+00
+ 6.51400e-08 0.00000e+00 6.51650e-08 6.70000e-04 6.52000e-08 0.00000e+00
+ 6.53400e-08 0.00000e+00 6.53650e-08 6.70000e-04 6.54000e-08 0.00000e+00
+ 6.55400e-08 0.00000e+00 6.55650e-08 6.70000e-04 6.56000e-08 0.00000e+00
+ 6.57400e-08 0.00000e+00 6.57650e-08 6.70000e-04 6.58000e-08 0.00000e+00
+ 6.59400e-08 0.00000e+00 6.59650e-08 6.70000e-04 6.60000e-08 0.00000e+00
+ 6.61400e-08 0.00000e+00 6.61650e-08 6.70000e-04 6.62000e-08 0.00000e+00
+ 6.63400e-08 0.00000e+00 6.63650e-08 6.70000e-04 6.64000e-08 0.00000e+00
+ 6.65400e-08 0.00000e+00 6.65650e-08 6.70000e-04 6.66000e-08 0.00000e+00
+ 6.67400e-08 0.00000e+00 6.67650e-08 6.70000e-04 6.68000e-08 0.00000e+00
+ 6.69400e-08 0.00000e+00 6.69650e-08 6.70000e-04 6.70000e-08 0.00000e+00
+ 6.71400e-08 0.00000e+00 6.71650e-08 6.70000e-04 6.72000e-08 0.00000e+00
+ 6.73400e-08 0.00000e+00 6.73650e-08 6.70000e-04 6.74000e-08 0.00000e+00
+ 6.75400e-08 0.00000e+00 6.75650e-08 6.70000e-04 6.76000e-08 0.00000e+00
+ 6.77400e-08 0.00000e+00 6.77650e-08 6.70000e-04 6.78000e-08 0.00000e+00
+ 6.79400e-08 0.00000e+00 6.79650e-08 6.70000e-04 6.80000e-08 0.00000e+00
+ 6.81400e-08 0.00000e+00 6.81650e-08 6.70000e-04 6.82000e-08 0.00000e+00
+ 6.83400e-08 0.00000e+00 6.83650e-08 6.70000e-04 6.84000e-08 0.00000e+00
+ 6.85400e-08 0.00000e+00 6.85650e-08 6.70000e-04 6.86000e-08 0.00000e+00
+ 6.87400e-08 0.00000e+00 6.87650e-08 6.70000e-04 6.88000e-08 0.00000e+00
+ 6.89400e-08 0.00000e+00 6.89650e-08 6.70000e-04 6.90000e-08 0.00000e+00
+ 6.91400e-08 0.00000e+00 6.91650e-08 6.70000e-04 6.92000e-08 0.00000e+00
+ 6.93400e-08 0.00000e+00 6.93650e-08 6.70000e-04 6.94000e-08 0.00000e+00
+ 6.95400e-08 0.00000e+00 6.95650e-08 6.70000e-04 6.96000e-08 0.00000e+00
+ 6.97400e-08 0.00000e+00 6.97650e-08 6.70000e-04 6.98000e-08 0.00000e+00
+ 6.99400e-08 0.00000e+00 6.99650e-08 6.70000e-04 7.00000e-08 0.00000e+00
+ 7.01400e-08 0.00000e+00 7.01650e-08 6.70000e-04 7.02000e-08 0.00000e+00
+ 7.03400e-08 0.00000e+00 7.03650e-08 6.70000e-04 7.04000e-08 0.00000e+00
+ 7.05400e-08 0.00000e+00 7.05650e-08 6.70000e-04 7.06000e-08 0.00000e+00
+ 7.07400e-08 0.00000e+00 7.07650e-08 6.70000e-04 7.08000e-08 0.00000e+00
+ 7.09400e-08 0.00000e+00 7.09650e-08 6.70000e-04 7.10000e-08 0.00000e+00
+ 7.11400e-08 0.00000e+00 7.11650e-08 6.70000e-04 7.12000e-08 0.00000e+00
+ 7.13400e-08 0.00000e+00 7.13650e-08 6.70000e-04 7.14000e-08 0.00000e+00
+ 7.15400e-08 0.00000e+00 7.15650e-08 6.70000e-04 7.16000e-08 0.00000e+00
+ 7.17400e-08 0.00000e+00 7.17650e-08 6.70000e-04 7.18000e-08 0.00000e+00
+ 7.19400e-08 0.00000e+00 7.19650e-08 6.70000e-04 7.20000e-08 0.00000e+00
+ 7.21400e-08 0.00000e+00 7.21650e-08 6.70000e-04 7.22000e-08 0.00000e+00
+ 7.23400e-08 0.00000e+00 7.23650e-08 6.70000e-04 7.24000e-08 0.00000e+00
+ 7.25400e-08 0.00000e+00 7.25650e-08 6.70000e-04 7.26000e-08 0.00000e+00
+ 7.27400e-08 0.00000e+00 7.27650e-08 6.70000e-04 7.28000e-08 0.00000e+00
+ 7.29400e-08 0.00000e+00 7.29650e-08 6.70000e-04 7.30000e-08 0.00000e+00
+ 7.31400e-08 0.00000e+00 7.31650e-08 6.70000e-04 7.32000e-08 0.00000e+00
+ 7.33400e-08 0.00000e+00 7.33650e-08 6.70000e-04 7.34000e-08 0.00000e+00
+ 7.35400e-08 0.00000e+00 7.35650e-08 6.70000e-04 7.36000e-08 0.00000e+00
+ 7.37400e-08 0.00000e+00 7.37650e-08 6.70000e-04 7.38000e-08 0.00000e+00
+ 7.39400e-08 0.00000e+00 7.39650e-08 6.70000e-04 7.40000e-08 0.00000e+00
+ 7.41400e-08 0.00000e+00 7.41650e-08 6.70000e-04 7.42000e-08 0.00000e+00
+ 7.43400e-08 0.00000e+00 7.43650e-08 6.70000e-04 7.44000e-08 0.00000e+00
+ 7.45400e-08 0.00000e+00 7.45650e-08 6.70000e-04 7.46000e-08 0.00000e+00
+ 7.47400e-08 0.00000e+00 7.47650e-08 6.70000e-04 7.48000e-08 0.00000e+00
+ 7.49400e-08 0.00000e+00 7.49650e-08 6.70000e-04 7.50000e-08 0.00000e+00
+ 7.51400e-08 0.00000e+00 7.51650e-08 6.70000e-04 7.52000e-08 0.00000e+00
+ 7.53400e-08 0.00000e+00 7.53650e-08 6.70000e-04 7.54000e-08 0.00000e+00
+ 7.55400e-08 0.00000e+00 7.55650e-08 6.70000e-04 7.56000e-08 0.00000e+00
+ 7.57400e-08 0.00000e+00 7.57650e-08 6.70000e-04 7.58000e-08 0.00000e+00
+ 7.59400e-08 0.00000e+00 7.59650e-08 6.70000e-04 7.60000e-08 0.00000e+00
+ 7.61400e-08 0.00000e+00 7.61650e-08 6.70000e-04 7.62000e-08 0.00000e+00
+ 7.63400e-08 0.00000e+00 7.63650e-08 6.70000e-04 7.64000e-08 0.00000e+00
+ 7.65400e-08 0.00000e+00 7.65650e-08 6.70000e-04 7.66000e-08 0.00000e+00
+ 7.67400e-08 0.00000e+00 7.67650e-08 6.70000e-04 7.68000e-08 0.00000e+00
+ 7.69400e-08 0.00000e+00 7.69650e-08 6.70000e-04 7.70000e-08 0.00000e+00
+ 7.71400e-08 0.00000e+00 7.71650e-08 6.70000e-04 7.72000e-08 0.00000e+00
+ 7.73400e-08 0.00000e+00 7.73650e-08 6.70000e-04 7.74000e-08 0.00000e+00
+ 7.75400e-08 0.00000e+00 7.75650e-08 6.70000e-04 7.76000e-08 0.00000e+00
+ 7.77400e-08 0.00000e+00 7.77650e-08 6.70000e-04 7.78000e-08 0.00000e+00
+ 7.79400e-08 0.00000e+00 7.79650e-08 6.70000e-04 7.80000e-08 0.00000e+00
+ 7.81400e-08 0.00000e+00 7.81650e-08 6.70000e-04 7.82000e-08 0.00000e+00
+ 7.83400e-08 0.00000e+00 7.83650e-08 6.70000e-04 7.84000e-08 0.00000e+00
+ 7.85400e-08 0.00000e+00 7.85650e-08 6.70000e-04 7.86000e-08 0.00000e+00
+ 7.87400e-08 0.00000e+00 7.87650e-08 6.70000e-04 7.88000e-08 0.00000e+00
+ 7.89400e-08 0.00000e+00 7.89650e-08 6.70000e-04 7.90000e-08 0.00000e+00
+ 7.91400e-08 0.00000e+00 7.91650e-08 6.70000e-04 7.92000e-08 0.00000e+00
+ 7.93400e-08 0.00000e+00 7.93650e-08 6.70000e-04 7.94000e-08 0.00000e+00
+ 7.95400e-08 0.00000e+00 7.95650e-08 6.70000e-04 7.96000e-08 0.00000e+00
+ 7.97400e-08 0.00000e+00 7.97650e-08 6.70000e-04 7.98000e-08 0.00000e+00
+ 7.99400e-08 0.00000e+00 7.99650e-08 6.70000e-04 8.00000e-08 0.00000e+00
+ 8.01400e-08 0.00000e+00 8.01650e-08 6.70000e-04 8.02000e-08 0.00000e+00
+ 8.03400e-08 0.00000e+00 8.03650e-08 6.70000e-04 8.04000e-08 0.00000e+00
+ 8.05400e-08 0.00000e+00 8.05650e-08 6.70000e-04 8.06000e-08 0.00000e+00
+ 8.07400e-08 0.00000e+00 8.07650e-08 6.70000e-04 8.08000e-08 0.00000e+00
+ 8.09400e-08 0.00000e+00 8.09650e-08 6.70000e-04 8.10000e-08 0.00000e+00
+ 8.11400e-08 0.00000e+00 8.11650e-08 6.70000e-04 8.12000e-08 0.00000e+00
+ 8.13400e-08 0.00000e+00 8.13650e-08 6.70000e-04 8.14000e-08 0.00000e+00
+ 8.15400e-08 0.00000e+00 8.15650e-08 6.70000e-04 8.16000e-08 0.00000e+00
+ 8.17400e-08 0.00000e+00 8.17650e-08 6.70000e-04 8.18000e-08 0.00000e+00
+ 8.19400e-08 0.00000e+00 8.19650e-08 6.70000e-04 8.20000e-08 0.00000e+00
+ 8.21400e-08 0.00000e+00 8.21650e-08 6.70000e-04 8.22000e-08 0.00000e+00
+ 8.23400e-08 0.00000e+00 8.23650e-08 6.70000e-04 8.24000e-08 0.00000e+00
+ 8.25400e-08 0.00000e+00 8.25650e-08 6.70000e-04 8.26000e-08 0.00000e+00
+ 8.27400e-08 0.00000e+00 8.27650e-08 6.70000e-04 8.28000e-08 0.00000e+00
+ 8.29400e-08 0.00000e+00 8.29650e-08 6.70000e-04 8.30000e-08 0.00000e+00
+ 8.31400e-08 0.00000e+00 8.31650e-08 6.70000e-04 8.32000e-08 0.00000e+00
+ 8.33400e-08 0.00000e+00 8.33650e-08 6.70000e-04 8.34000e-08 0.00000e+00
+ 8.35400e-08 0.00000e+00 8.35650e-08 6.70000e-04 8.36000e-08 0.00000e+00
+ 8.37400e-08 0.00000e+00 8.37650e-08 6.70000e-04 8.38000e-08 0.00000e+00
+ 8.39400e-08 0.00000e+00 8.39650e-08 6.70000e-04 8.40000e-08 0.00000e+00
+ 8.41400e-08 0.00000e+00 8.41650e-08 6.70000e-04 8.42000e-08 0.00000e+00
+ 8.43400e-08 0.00000e+00 8.43650e-08 6.70000e-04 8.44000e-08 0.00000e+00
+ 8.45400e-08 0.00000e+00 8.45650e-08 6.70000e-04 8.46000e-08 0.00000e+00
+ 8.47400e-08 0.00000e+00 8.47650e-08 6.70000e-04 8.48000e-08 0.00000e+00
+ 8.49400e-08 0.00000e+00 8.49650e-08 6.70000e-04 8.50000e-08 0.00000e+00
+ 8.51400e-08 0.00000e+00 8.51650e-08 6.70000e-04 8.52000e-08 0.00000e+00
+ 8.53400e-08 0.00000e+00 8.53650e-08 6.70000e-04 8.54000e-08 0.00000e+00
+ 8.55400e-08 0.00000e+00 8.55650e-08 6.70000e-04 8.56000e-08 0.00000e+00
+ 8.57400e-08 0.00000e+00 8.57650e-08 6.70000e-04 8.58000e-08 0.00000e+00
+ 8.59400e-08 0.00000e+00 8.59650e-08 6.70000e-04 8.60000e-08 0.00000e+00
+ 8.61400e-08 0.00000e+00 8.61650e-08 6.70000e-04 8.62000e-08 0.00000e+00
+ 8.63400e-08 0.00000e+00 8.63650e-08 6.70000e-04 8.64000e-08 0.00000e+00
+ 8.65400e-08 0.00000e+00 8.65650e-08 6.70000e-04 8.66000e-08 0.00000e+00
+ 8.67400e-08 0.00000e+00 8.67650e-08 6.70000e-04 8.68000e-08 0.00000e+00
+ 8.69400e-08 0.00000e+00 8.69650e-08 6.70000e-04 8.70000e-08 0.00000e+00
+ 8.71400e-08 0.00000e+00 8.71650e-08 6.70000e-04 8.72000e-08 0.00000e+00
+ 8.73400e-08 0.00000e+00 8.73650e-08 6.70000e-04 8.74000e-08 0.00000e+00
+ 8.75400e-08 0.00000e+00 8.75650e-08 6.70000e-04 8.76000e-08 0.00000e+00
+ 8.77400e-08 0.00000e+00 8.77650e-08 6.70000e-04 8.78000e-08 0.00000e+00
+ 8.79400e-08 0.00000e+00 8.79650e-08 6.70000e-04 8.80000e-08 0.00000e+00
+ 8.81400e-08 0.00000e+00 8.81650e-08 6.70000e-04 8.82000e-08 0.00000e+00
+ 8.83400e-08 0.00000e+00 8.83650e-08 6.70000e-04 8.84000e-08 0.00000e+00
+ 8.85400e-08 0.00000e+00 8.85650e-08 6.70000e-04 8.86000e-08 0.00000e+00
+ 8.87400e-08 0.00000e+00 8.87650e-08 6.70000e-04 8.88000e-08 0.00000e+00
+ 8.89400e-08 0.00000e+00 8.89650e-08 6.70000e-04 8.90000e-08 0.00000e+00
+ 8.91400e-08 0.00000e+00 8.91650e-08 6.70000e-04 8.92000e-08 0.00000e+00
+ 8.93400e-08 0.00000e+00 8.93650e-08 6.70000e-04 8.94000e-08 0.00000e+00
+ 8.95400e-08 0.00000e+00 8.95650e-08 6.70000e-04 8.96000e-08 0.00000e+00
+ 8.97400e-08 0.00000e+00 8.97650e-08 6.70000e-04 8.98000e-08 0.00000e+00
+ 8.99400e-08 0.00000e+00 8.99650e-08 6.70000e-04 9.00000e-08 0.00000e+00
+ 9.01400e-08 0.00000e+00 9.01650e-08 6.70000e-04 9.02000e-08 0.00000e+00
+ 9.03400e-08 0.00000e+00 9.03650e-08 6.70000e-04 9.04000e-08 0.00000e+00
+ 9.05400e-08 0.00000e+00 9.05650e-08 6.70000e-04 9.06000e-08 0.00000e+00
+ 9.07400e-08 0.00000e+00 9.07650e-08 6.70000e-04 9.08000e-08 0.00000e+00
+ 9.09400e-08 0.00000e+00 9.09650e-08 6.70000e-04 9.10000e-08 0.00000e+00
+ 9.11400e-08 0.00000e+00 9.11650e-08 6.70000e-04 9.12000e-08 0.00000e+00
+ 9.13400e-08 0.00000e+00 9.13650e-08 6.70000e-04 9.14000e-08 0.00000e+00
+ 9.15400e-08 0.00000e+00 9.15650e-08 6.70000e-04 9.16000e-08 0.00000e+00
+ 9.17400e-08 0.00000e+00 9.17650e-08 6.70000e-04 9.18000e-08 0.00000e+00
+ 9.19400e-08 0.00000e+00 9.19650e-08 6.70000e-04 9.20000e-08 0.00000e+00
+ 9.21400e-08 0.00000e+00 9.21650e-08 6.70000e-04 9.22000e-08 0.00000e+00
+ 9.23400e-08 0.00000e+00 9.23650e-08 6.70000e-04 9.24000e-08 0.00000e+00
+ 9.25400e-08 0.00000e+00 9.25650e-08 6.70000e-04 9.26000e-08 0.00000e+00
+ 9.27400e-08 0.00000e+00 9.27650e-08 6.70000e-04 9.28000e-08 0.00000e+00
+ 9.29400e-08 0.00000e+00 9.29650e-08 6.70000e-04 9.30000e-08 0.00000e+00
+ 9.31400e-08 0.00000e+00 9.31650e-08 6.70000e-04 9.32000e-08 0.00000e+00
+ 9.33400e-08 0.00000e+00 9.33650e-08 6.70000e-04 9.34000e-08 0.00000e+00
+ 9.35400e-08 0.00000e+00 9.35650e-08 6.70000e-04 9.36000e-08 0.00000e+00
+ 9.37400e-08 0.00000e+00 9.37650e-08 6.70000e-04 9.38000e-08 0.00000e+00
+ 9.39400e-08 0.00000e+00 9.39650e-08 6.70000e-04 9.40000e-08 0.00000e+00
+ 9.41400e-08 0.00000e+00 9.41650e-08 6.70000e-04 9.42000e-08 0.00000e+00
+ 9.43400e-08 0.00000e+00 9.43650e-08 6.70000e-04 9.44000e-08 0.00000e+00
+ 9.45400e-08 0.00000e+00 9.45650e-08 6.70000e-04 9.46000e-08 0.00000e+00
+ 9.47400e-08 0.00000e+00 9.47650e-08 6.70000e-04 9.48000e-08 0.00000e+00
+ 9.49400e-08 0.00000e+00 9.49650e-08 6.70000e-04 9.50000e-08 0.00000e+00
+ 9.51400e-08 0.00000e+00 9.51650e-08 6.70000e-04 9.52000e-08 0.00000e+00
+ 9.53400e-08 0.00000e+00 9.53650e-08 6.70000e-04 9.54000e-08 0.00000e+00
+ 9.55400e-08 0.00000e+00 9.55650e-08 6.70000e-04 9.56000e-08 0.00000e+00
+ 9.57400e-08 0.00000e+00 9.57650e-08 6.70000e-04 9.58000e-08 0.00000e+00
+ 9.59400e-08 0.00000e+00 9.59650e-08 6.70000e-04 9.60000e-08 0.00000e+00
+ 9.61400e-08 0.00000e+00 9.61650e-08 6.70000e-04 9.62000e-08 0.00000e+00
+ 9.63400e-08 0.00000e+00 9.63650e-08 6.70000e-04 9.64000e-08 0.00000e+00
+ 9.65400e-08 0.00000e+00 9.65650e-08 6.70000e-04 9.66000e-08 0.00000e+00
+ 9.67400e-08 0.00000e+00 9.67650e-08 6.70000e-04 9.68000e-08 0.00000e+00
+ 9.69400e-08 0.00000e+00 9.69650e-08 6.70000e-04 9.70000e-08 0.00000e+00
+ 9.71400e-08 0.00000e+00 9.71650e-08 6.70000e-04 9.72000e-08 0.00000e+00
+ 9.73400e-08 0.00000e+00 9.73650e-08 6.70000e-04 9.74000e-08 0.00000e+00
+ 9.75400e-08 0.00000e+00 9.75650e-08 6.70000e-04 9.76000e-08 0.00000e+00
+ 9.77400e-08 0.00000e+00 9.77650e-08 6.70000e-04 9.78000e-08 0.00000e+00
+ 9.79400e-08 0.00000e+00 9.79650e-08 6.70000e-04 9.80000e-08 0.00000e+00
+ 9.81400e-08 0.00000e+00 9.81650e-08 6.70000e-04 9.82000e-08 0.00000e+00
+ 9.83400e-08 0.00000e+00 9.83650e-08 6.70000e-04 9.84000e-08 0.00000e+00
+ 9.85400e-08 0.00000e+00 9.85650e-08 6.70000e-04 9.86000e-08 0.00000e+00
+ 9.87400e-08 0.00000e+00 9.87650e-08 6.70000e-04 9.88000e-08 0.00000e+00
+ 9.89400e-08 0.00000e+00 9.89650e-08 6.70000e-04 9.90000e-08 0.00000e+00
+ 9.91400e-08 0.00000e+00 9.91650e-08 6.70000e-04 9.92000e-08 0.00000e+00
+ 9.93400e-08 0.00000e+00 9.93650e-08 6.70000e-04 9.94000e-08 0.00000e+00
+ 9.95400e-08 0.00000e+00 9.95650e-08 6.70000e-04 9.96000e-08 0.00000e+00
+ 9.97400e-08 0.00000e+00 9.97650e-08 6.70000e-04 9.98000e-08 0.00000e+00
+ 9.99400e-08 0.00000e+00 9.99650e-08 6.70000e-04 1.00000e-07 0.00000e+00
+ 1.00140e-07 0.00000e+00 1.00165e-07 6.70000e-04 1.00200e-07 0.00000e+00
+ 1.00340e-07 0.00000e+00 1.00365e-07 6.70000e-04 1.00400e-07 0.00000e+00
+ 1.00540e-07 0.00000e+00 1.00565e-07 6.70000e-04 1.00600e-07 0.00000e+00)

.subckt SYNAPSEfastestnext2 DIN DOUTL DOUTR WEIGHTL WEIGHTR NODEM 
LINPUT DIN 0 5.25p
#RINPUT DINX 0 0.5

LSTORE1 WEIGHTL NODEM 45.8p
LSTORE2 NODEM WEIGHTR 45.8p
KWEIGHT1 LWIN LSTORE1  -0.1
#KWEIGHT1 LWIN LSTORE1  -0.05
LWin 0 MIDDLE  40p
L1 LEFT MIDDLE 5p
L2 MIDDLE RIGHT 5p
.param shunt = 6
RSHUNT1 LEFT 0 shunt
RSHUNT2 RIGHT 0 shunt
#WAS 5.3
B1 LEFT 3par N1 jjmit area=0.5
B2 RIGHT 4par N2 jjmit area=0.5
LP1 3par 0 0.2p
LP2 4par 0 0.2p
LQ MIDDLE 0 20.84p
#LQ MIDDLE 0 40.84p
K1 L2  LINPUT -0.25
K2 LINPUT L1 -0.25
KOUT LQ LOUT -0.01
#WAS 35
LOUT DOUTL DOUTR 25P
#consider taking out lout but how do I couple then...
.ends SYNAPSEfastestnext2
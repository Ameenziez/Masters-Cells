.SUBCKT NEURONLETTER INPUT1 INPUT2 INPUT3 INPUT4 INPUT5 INPUT6 INPUT7 INPUT8 INPUT9 INPUTB TARGET INITIAL1 INITIAL2 INITIAL3 INITIAL4 INITIAL5 INITIAL6 INITIAL7 INITIAL8 INITIAL9 INITIALB XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT DCCONVIN DCCONVOUT  CONSTIN
#took out DOUTCOMP
Lin1 INPUT1 IN12 10p
LINFeed1 0 INADJUST1 10p
Kin1 LIN1 LINFeed1 -0.01

Lin2 INPUT2 IN22 10p
LINFeed2 0 INADJUST2 10p
Kin2 LIN2 LINFeed2 -0.01

Lin3 INPUT3 IN32 10p
LINFeed3 0 INADJUST3 10p
Kin3 LIN3 LINFeed3 -0.01

Lin4 INPUT4 IN42 10p
LINFeed4 0 INADJUST4 10p
Kin4 LIN4 LINFeed4 -0.01

Lin5 INPUT5 IN52 10p
LINFeed5 0 INADJUST5 10p
Kin5 LIN5 LINFeed5 -0.01

Lin6 INPUT6 IN62 10p
LINFeed6 0 INADJUST6 10p
Kin6 LIN6 LINFeed6 -0.01

Lin7 INPUT7 IN72 10p
LINFeed7 0 INADJUST7 10p
Kin7 LIN7 LINFeed7 -0.01

Lin8 INPUT8 IN82 10p
LINFeed8 0 INADJUST8 10p
Kin8 LIN8 LINFeed8 -0.01

Lin9 INPUT9 IN92 10p
LINFeed9 0 INADJUST9 10p
Kin9 LIN9 LINFeed9 -0.01



Ltarget TARGET 0 10p
LtargetFeed1 0 TARGETIN1 10p
LtargetFeed2 0 TARGETIN2 10p
LtargetFeed3 0 TARGETIN3 10p
LtargetFeed4 0 TARGETIN4 10p
LtargetFeed5 0 TARGETIN5 10p
LtargetFeed6 0 TARGETIN6 10p
LtargetFeed7 0 TARGETIN7 10p
LtargetFeed8 0 TARGETIN8 10p
LtargetFeed9 0 TARGETIN9 10p
LtargetFeed10 0 TARGETINB 10p
Ktarget1 Ltarget LtargetFeed1 -0.01
Ktarget2 Ltarget LtargetFeed2 -0.01
Ktarget3 Ltarget LtargetFeed3 -0.01
Ktarget4 Ltarget LtargetFeed4 -0.01
Ktarget5 Ltarget LtargetFeed5 -0.01
Ktarget6 Ltarget LtargetFeed6 -0.01
Ktarget7 Ltarget LtargetFeed7 -0.01
Ktarget8 Ltarget LtargetFeed8 -0.01
Ktarget9 Ltarget LtargetFeed9 -0.01
Ktarget10 Ltarget LtargetFeed10 -0.01


LinBIAS INPUTB INB2 10p
LINBIASFEED 0 INADJUSTBIAS 10p
KinBIAS1 LINBIAS LINBIASFeed -0.01


XSYN1 SYNAPSEfastest IN12 OUTL1 OUTL2 WEIGHTL1 WEIGHTR1 INITIAL1
XSTORE1 BISTORE WPLUS1 WMINUS1 WEIGHTL1 WEIGHTR1
XSYN2 SYNAPSEfastest IN22 OUTL2 OUTL3 WEIGHTL2 WEIGHTR2 INITIAL2
XSTORE2 BISTORE WPLUS2 WMINUS2 WEIGHTL2 WEIGHTR2
XSYN3 SYNAPSEfastest IN32 OUTL3 OUTL4 WEIGHTL3 WEIGHTR3 INITIAL3
XSTORE3 BISTORE WPLUS3 WMINUS3 WEIGHTL3 WEIGHTR3
XSYN4 SYNAPSEfastest IN42 OUTL4 OUTL5 WEIGHTL4 WEIGHTR4 INITIAL4
XSTORE4 BISTORE WPLUS4 WMINUS4 WEIGHTL4 WEIGHTR4
XSYN5 SYNAPSEfastest IN52 OUTL5 OUTL6 WEIGHTL5 WEIGHTR5 INITIAL5
XSTORE5 BISTORE WPLUS5 WMINUS5 WEIGHTL5 WEIGHTR5
XSYN6 SYNAPSEfastest IN62 OUTL6 OUTL7 WEIGHTL6 WEIGHTR6 INITIAL6
XSTORE6 BISTORE WPLUS6 WMINUS6 WEIGHTL6 WEIGHTR6
XSYN7 SYNAPSEfastest IN72 OUTL7 OUTL8 WEIGHTL7 WEIGHTR7 INITIAL7
XSTORE7 BISTORE WPLUS7 WMINUS7 WEIGHTL7 WEIGHTR7
XSYN8 SYNAPSEfastest IN82 OUTL8 OUTL9 WEIGHTL8 WEIGHTR8 INITIAL8
XSTORE8 BISTORE WPLUS8 WMINUS8 WEIGHTL8 WEIGHTR8
XSYN9 SYNAPSEfastest IN92 OUTL9 OUTL10 WEIGHTL9 WEIGHTR9 INITIAL9
XSTORE9 BISTORE WPLUS9 WMINUS9 WEIGHTL9 WEIGHTR9
XSYNBIAS SYNAPSEfastest INB2 OUTL10 0 WEIGHTLB WEIGHTRB INITIALB
XSTOREBIAS BISTORE WPLUSB WMINUSB WEIGHTLB WEIGHTRB

#ACTIVATION
#XCOMP COMP20 XIN1 OUTL1 A4 DCIN DC4 0 DOUTCOMP 0 ADJUSTBACK1P 0 0 ADJUSTBACK1N ADJUSTBACK2P 0 0 ADJUSTBACK2N ADJUSTBACK3P 0 0 ADJUSTBACK3N  ADJUSTBACK4P 0 0 ADJUSTBACK4N  ADJUSTBACK5P 0 0 ADJUSTBACK5N  ADJUSTBACK6P 0 0 ADJUSTBACK6N  ADJUSTBACK7P 0 0 ADJUSTBACK7N  ADJUSTBACK8P 0 0 ADJUSTBACK8N ADJUSTBACK9P 0 0 ADJUSTBACK9N  ADJUSTBIASP 0  0 ADJUSTBIASN  CONSTIN
XCOMP COMP20 XIN1 OUTL1 A4 DCIN DC4  ADJUSTBACK1N 0  0 ADJUSTBACK1P ADJUSTBACK2N 0 0 ADJUSTBACK2P ADJUSTBACK3N 0 0 ADJUSTBACK3P  ADJUSTBACK4N 0 0 ADJUSTBACK4P  ADJUSTBACK5N 0 0 ADJUSTBACK5P  ADJUSTBACK6N 0 0 ADJUSTBACK6P  ADJUSTBACK7N 0 0 ADJUSTBACK7P  ADJUSTBACK8N 0 0 ADJUSTBACK8P ADJUSTBACK9N 0 0 ADJUSTBACK9P  ADJUSTBACKBIASN 0  0 ADJUSTBACKBIASP  CONSTIN


#need to reverse some polarities... does't seem to be able to decrement
# WEIGHT ADJUSTMENT

#XADJUST1 ADJUSTNEW2 A4 A5 XIN2 B4 INADJUST1 ADJUSTBACK1 TARGETIN1    DC4 DC5     INCR1 DECR1
#XADJUST2 ADJUSTNEW2 A5 A6  B4 B5  INADJUST2 ADJUSTBACK2 TARGETIN2  DC5 DC6     INCR2 DECR2
#XADJUSTB ADJUSTNEW2 A6 A7  B5 B6  INADJUSTBIAS ADJUSTBIAS TARGETINB DC6  DC7      INCRB DECRB
#XADJUST3 ADJUSTNEW2 A7 A8 B6 B7 INADJUST3 ADJUSTBACK3 TARGETIN3    DC7 DC8     INCR3 DECR3
#XADJUST4 ADJUSTNEW2 A8 A9  B7 B8  INADJUST4 ADJUSTBACK4 TARGETIN4  DC8 DC9     INCR4 DECR4
#XADJUST5 ADJUSTNEW2 A9 A10  B8 B9  INADJUST5 ADJUSTBACK5 TARGETIN5 DC9  DC10      INCR5 DECR5
#XADJUST6 ADJUSTNEW2 A10 A11 B9 B10 INADJUST6 ADJUSTBACK6 TARGETIN6    DC10 DC11     INCR6 DECR6
#XADJUST7 ADJUSTNEW2 A11 A12  B10 B11  INADJUST7 ADJUSTBACK7 TARGETIN7  DC11 DC12     INCR7 DECR7
#XADJUST8 ADJUSTNEW2 A12 A13  B11 B12  INADJUST8 ADJUSTBACK8 TARGETIN8 DC12  DC13      INCR8 DECR8
#XADJUST9 ADJUSTNEW2 A13 XOUT1  B12 B13  INADJUST9 ADJUSTBACK9 TARGETIN9 DC13  DCOUT      INCR9 DECR9

#REVERSED DCS HERE
#XPERCEPTRON11 PERCEPTRON  A4 A5  XIN2 B1  INADJUST1 ADJUSTBACK1P ADJUSTBACK1N TARGETIN1 DC5 DC4 DECR1 INCR1 
#XPERCEPTRON12 PERCEPTRON  A5 A6  B1 B2  INADJUST2 ADJUSTBACK2P ADJUSTBACK2N  TARGETIN2 DC6 DC5  DECR2 INCR2
#XPERCEPTRON13 PERCEPTRON  A6 A7  B2 B3  INADJUST3 ADJUSTBACK3P ADJUSTBACK3N  TARGETIN3 DC7 DC6  DECR3 INCR3
#XPERCEPTRON14 PERCEPTRON  A7 A8  B3 B4  INADJUST4 ADJUSTBACK4P ADJUSTBACK4N  TARGETIN4 DC8 DC7  DECR4 INCR4
#XPERCEPTRON15 PERCEPTRON  A8 A9  B4 B5  INADJUST5 ADJUSTBACK5P ADJUSTBACK5N  TARGETIN5 DC9 DC8  DECR5 INCR5
#XPERCEPTRON16 PERCEPTRON  A9 A10  B5 B6  INADJUST6 ADJUSTBACK6P ADJUSTBACK6N  TARGETIN6 DC10 DC9  DECR6 INCR6
#XPERCEPTRON17 PERCEPTRON  A10 A11  B6 B7  INADJUST7 ADJUSTBACK7P ADJUSTBACK7N  TARGETIN7 DC11 DC10  DECR7 INCR7
#XPERCEPTRON18 PERCEPTRON  A11 A12  B7 B8  INADJUST8 ADJUSTBACK8P ADJUSTBACK8N  TARGETIN8 DC12 DC11  DECR8 INCR8
#XPERCEPTRON19 PERCEPTRON  A12 A13  B8 B9  INADJUST9 ADJUSTBACK9P ADJUSTBACK9N  TARGETIN9 DC13 DC12  DECR9 INCR9
#XPERCEPTRONB PERCEPTRON  A13 XOUT1  B9 B10  INADJUSTBIAS ADJUSTBACKBIASP ADJUSTBACKBIASN  TARGETINB  DCOUT DC13   DECRB INCRB

XPERCEPTRON11 PERCEPTRON3  A4 A5  XIN2 B1  INADJUST1 ADJUSTBACK1N ADJUSTBACK1P TARGETIN1 DC5 DC4 INCR1 DECR1 
XPERCEPTRON12 PERCEPTRON3  A5 A6  B1 B2  INADJUST2 ADJUSTBACK2N ADJUSTBACK2P  TARGETIN2 DC6 DC5  INCR2 DECR2
XPERCEPTRON13 PERCEPTRON3  A6 A7  B2 B3  INADJUST3 ADJUSTBACK3N ADJUSTBACK3P  TARGETIN3 DC7 DC6  INCR3 DECR3
XPERCEPTRON14 PERCEPTRON3  A7 A8  B3 B4  INADJUST4 ADJUSTBACK4N ADJUSTBACK4P  TARGETIN4 DC8 DC7  INCR4 DECR4
XPERCEPTRON15 PERCEPTRON3  A8 A9  B4 B5  INADJUST5 ADJUSTBACK5N ADJUSTBACK5P  TARGETIN5 DC9 DC8  INCR5 DECR5
XPERCEPTRON16 PERCEPTRON3  A9 A10  B5 B6  INADJUST6 ADJUSTBACK6N ADJUSTBACK6P  TARGETIN6 DC10 DC9  INCR6 DECR6
XPERCEPTRON17 PERCEPTRON3  A10 A11  B6 B7  INADJUST7 ADJUSTBACK7N ADJUSTBACK7P  TARGETIN7 DC11 DC10  INCR7 DECR7
XPERCEPTRON18 PERCEPTRON3  A11 A12  B7 B8  INADJUST8 ADJUSTBACK8N ADJUSTBACK8P  TARGETIN8 DC12 DC11  INCR8 DECR8
XPERCEPTRON19 PERCEPTRON3  A12 A13  B8 B9  INADJUST9 ADJUSTBACK9N ADJUSTBACK9P  TARGETIN9 DC13 DC12  INCR9 DECR9
XPERCEPTRONB PERCEPTRON3  A13 XOUT1  B9 B10  INADJUSTBIAS ADJUSTBACKBIASN ADJUSTBACKBIASP  TARGETINB  DCOUT DC13   INCRB DECRB



#XCONV1 CONV B13 B14 DCC4 DCCONVIN     INCR1 DECR1 WPLUS1 WMINUS1
#XCONV2 CONV B14 B15 DCc5 DCc4         INCR2 DECR2 WPLUS2 WMINUS2
#XCONVB CONV B15 B16 DCC6 DCc5         INCRB DECRB WPLUSB WMINUSB
#XCONV3 CONV B16 B17 DCC7 DCC6         INCR3 DECR3 WPLUS3 WMINUS3
#XCONV4 CONV B17 B18 DCc8 DCc7         INCR4 DECR4 WPLUS4 WMINUS4
#XCONV5 CONV B18 B19 DCC9 DCC8         INCR5 DECR5 WPLUS5 WMINUS5
#XCONV6 CONV B19 B20 DCc10 DCc9        INCR6 DECR6 WPLUS6 WMINUS6
#XCONV7 CONV B20 B21 DCC11 DCC10       INCR7 DECR7 WPLUS7 WMINUS7
#XCONV8 CONV B21 B22 DCc12 DCc11       INCR8 DECR8 WPLUS8 WMINUS8
#XCONV9 CONV B22 XOUT2 DCCONVOUT DCc12 INCR9 DECR9 WPLUS9 WMINUS9

#XCONV1 CONV A15 A14  DCC4  DCCONVIN     INCR1 DECR1 WPLUS1 WMINUS1
#XCONV2 CONV A16 A15 DCc5 DCc4         INCR2 DECR2 WPLUS2 WMINUS2
#XCONVB CONV A17 A16  DCC6 DCc5         INCRB DECRB WPLUSB WMINUSB
#XCONV3 CONV A18 A17  DCC7 DCC6         INCR3 DECR3 WPLUS3 WMINUS3
#XCONV4 CONV A19 A18  DCc8 DCc7         INCR4 DECR4 WPLUS4 WMINUS4
#XCONV5 CONV A20 A19  DCC9 DCC8         INCR5 DECR5 WPLUS5 WMINUS5
#XCONV6 CONV A21 A20  DCc10 DCc9        INCR6 DECR6 WPLUS6 WMINUS6
#XCONV7 CONV A22 A21  DCC11 DCC10       INCR7 DECR7 WPLUS7 WMINUS7
#XCONV8 CONV A23 A22   DCc12 DCc11       INCR8 DECR8 WPLUS8 WMINUS8
#XCONV9 CONV XOUT1 A23  DCCONVOUT DCc12 INCR9 DECR9 WPLUS9 WMINUS9

XCONV1 CONV  B10 B11  DCC4 DCCONVIN    INCR1 DECR1 WPLUS1 WMINUS1
XCONV2 CONV B11 B12 DCc5 DCc4         INCR2 DECR2 WPLUS2 WMINUS2
XCONVB CONV B12 B13  DCC6 DCc5         INCRB DECRB WPLUSB WMINUSB
XCONV3 CONV B13 B14  DCC7 DCC6         INCR3 DECR3 WPLUS3 WMINUS3
XCONV4 CONV B14 B15  DCc8 DCc7         INCR4 DECR4 WPLUS4 WMINUS4
XCONV5 CONV B15 B16  DCC9 DCC8         INCR5 DECR5 WPLUS5 WMINUS5
XCONV6 CONV B16 B17  DCc10 DCc9        INCR6 DECR6 WPLUS6 WMINUS6
XCONV7 CONV B17 B18  DCC11 DCC10       INCR7 DECR7 WPLUS7 WMINUS7
XCONV8 CONV B18 B19   DCc12 DCc11       INCR8 DECR8 WPLUS8 WMINUS8
XCONV9 CONV B19 XOUT2  DCCONVOUT DCc12 INCR9 DECR9 WPLUS9 WMINUS9

.ENDS NEURONLETTER


.subckt COMP20 XIN DIN XOUT DCIN DCOUT DOUTL1 DOUTR1 DOUTL2 DOUTR2 DOUTL3 DOUTR3 DOUTL4 DOUTR4 DOUTL5 DOUTR5 DOUTL6 DOUTR6 DOUTL7 DOUTR7 DOUTL8 DOUTR8 DOUTL9 DOUTR9 DOUTL10 DOUTR10 DOUTL11 DOUTR11 DOUTL12 DOUTR12 DOUTL13 DOUTR13 DOUTL14 DOUTR14 DOUTL15 DOUTR15 DOUTL16 DOUTR16 DOUTL17 DOUTR17 DOUTL18 DOUTR18 DOUTL19 DOUTR19 DOUTL20 DOUTR20 CONSTIN
#iconst 0 CONST PWL(0 0 20p 47u)
#45 WORKS CURRENT CONFIG and or nor but nand a little sus, 47 WORKS ALL
Lconst CONSTIN 0 20p
#WAS CONSTIN
Lconstout 7Q 7 25.5P
Kconst  Lconst Lconstout 0.1
B1 8 0 11 jjmit area=0.5
B2 9 0 12 jjmit area=0.5
K1 LX LD 0.1322
K2 LD LOUT1 3.27E-5
K3 LX LOUT1 3.68E-5
K4 LD LQ 4.9E-4
K5 LX LQ 5.11E-4
K6 LOUT1 LQ 0.05
K7 L2 LD -0.1556
K8 L2 LX -0.228
K9 LX L1 -0.2284
K10 LD L1 -0.15559
K11 LD LOUT2 3.27E-5
K12 LX LOUT2 3.68E-5
K13 LOUT2 LQ 0.05
K14 LD LOUT3 3.27E-5
K15 LX LOUT3 3.68E-5
K16 LOUT3 LQ 0.05
K17 LD LOUT4 3.27E-5
K18 LX LOUT4 3.68E-5
K19 LOUT4 LQ 0.05
K20 LD LOUT5 3.27E-5
K21 LX LOUT5 3.68E-5
K22 LOUT5 LQ 0.05
K23 LD LOUT6 3.27E-5
K24 LX LOUT6 3.68E-5
K25 LOUT6 LQ 0.05
K26 LD LOUT7 3.27E-5
K27 LX LOUT7 3.68E-5
K28 LOUT7 LQ 0.05
K29 LD LOUT8 3.27E-5
K30 LX LOUT8 3.68E-5
K31 LOUT8 LQ 0.05
K29 LD LOUT9 3.27E-5
K30 LX LOUT9 3.68E-5
K31 LOUT9 LQ 0.05
K32 LD LOUT10 3.27E-5
K33 LX LOUT10 3.68E-5
K34 LOUT10 LQ 0.05
K35 LD LOUT11 3.27E-5
K36 LX LOUT11 3.68E-5
K37 LOUT11 LQ 0.05
K40 LOUT12 LQ 0.05
K41 LD LOUT12 3.27E-5
K42 LX LOUT12 3.68E-5
K43 LOUT13 LQ 0.05
K44 LD LOUT13 3.27E-5
K45 LX LOUT13 3.68E-5
K46 LOUT14 LQ 0.05
K47 LD LOUT14 3.27E-5
K48 LX LOUT14 3.68E-5
K49 LOUT15 LQ 0.05
K50 LD LOUT15 3.27E-5
K51 LX LOUT15 3.68E-5
K52 LOUT16 LQ 0.05
K53 LD LOUT16 3.27E-5
K54 LX LOUT16 3.68E-5
K55 LOUT17 LQ 0.05
K56 LD LOUT17 3.27E-5
K57 LX LOUT17 3.68E-5
K58 LOUT18 LQ 0.05
K59 LD LOUT18 3.27E-5
K60 LX LOUT18 3.68E-5
K61 LD LOUT19 3.27E-5
K62 LX LOUT19 3.68E-5
K63 LOUT19 LQ 0.05
K64 LD LOUT20 3.27E-5
K65 LX LOUT20 3.68E-5
K66 LOUT20 LQ 0.05

L1 8 7 1.51p
L2 7 9 1.51p
#LD DCIN DCOUT 7.94p
LD DCIN DCOUT 7.94p
LIN DIN 7Q 1.526p


#RSHUNT2 9 0 6
#WAS 6

LOUT1 DOUTL1 DOUTR1 20p
LOUT2 DOUTL2 DOUTR2 20P
LOUT3 DOUTL3 DOUTR3 20P
LOUT4 DOUTL4 DOUTR4 20P
LOUT5 DOUTL5 DOUTR5 20p
LOUT6 DOUTL6 DOUTR6 20P
LOUT7 DOUTL7 DOUTR7 20P
LOUT8 DOUTL8 DOUTR8 20P
LOUT9 DOUTL9 DOUTR9 20P
LOUT10 DOUTL10 DOUTR10 20P
LOUT11 DOUTL11 DOUTR11 20P
LOUT12 DOUTL12 DOUTR12 20P
LOUT13 DOUTL13 DOUTR13 20P
LOUT14 DOUTL14 DOUTR14 20P
LOUT15 DOUTL15 DOUTR15 20P
LOUT16 DOUTL16 DOUTR16 20P
LOUT17 DOUTL17 DOUTR17 20P
LOUT18 DOUTL18 DOUTR18 20P
LOUT19 DOUTL19 DOUTR19 20P
LOUT20 DOUTL20 DOUTR20 20P
LQ 7 0 28.84p
#WAS 5.84
LX XIN XOUT 6.51p
#LX XIN XOUT 9.51p
.ends COMP20

#works well!
#got the data to propagate
.include LSmitll_DCSFQ_PTLTX_v1p5.cir
.include LSmitll_bufft_v1p5.cir
.include LSmitll_PTLRX_SFQDC_v1p5.cir
.include LSmitll_SPLITT_v1p5.cir
.INCLUDE LSMITLL_JTLT_V1P5.CIR
.INCLUDE LSMITLL_MERGET_V1P5.CIR
.include storeedit.cir
.INCLUDE COMPONENTSEDIT.CIR
.INCLUDE COMP3.CIR
.INCLUDE COMP4.CIR
.INCLUDE COMP5.CIR
.INCLUDE COMP6.CIR
.include conv.cir
.INCLUDE synapsenext2.CIR
.INCLUDE DCPULSER.CIR
.INCLUDE MULTISPLIT.CIR
.include transmit.cir
.INCLUDE DELAY7.CIR
.INCLUDE AND.CIR
.INCLUDE AND3.CIR
.INCLUDE OR3.CIR
.include PERCEPTRON.CIR
.include CONVINTERFACE.cir


# TRY SHIFTING CLK OF OUTPUT BACK A BIT...

.tran 1ps 15000PS 0ps 1p
#MLP:
#D=Oi.T + Oi.!Oj + T.!Oj 

#setup circuitry
VAC1   A1   0   SIN(0 723mV 10GHz 200Ps 0)
RAC1   A1   A2   1000
LAC1   A2   A3   0.1p
VAC2   B1   0   SIN(0 723mV 10GHz 175.0ps 0)
RAC2   B1   B2   1000
LAC2   B2   B3   0.1p
VDC    DC1   0   pwl(0 0 20p 1023mV)
RDC    DC1   DC2   1000
LDC    DC2   DC3  0.1p
VDCconv    DCc1   0   PWL(0ps 0mV 20ps 1023mV 1.881e-08 1023mV 1.8811000000000002e-08 0)
RDCconv    DCc1   DCc2  640
LDCconv    DCc2   DCc3   0.1p




#SECOND LAYER SYNAPSE 1
IINITAL21 0 INITIAL21 PWL( 0 0 20P 0*2*22.6U)
XSTORE21 BISTORE SFQOUTPLUS21 SFQOUTMINUS21 WEIGHTL21 WEIGHTR21


#NEXT LAYER BIAS
#Iactualsynbias21 0 ACTUALSYNB21x PWL(0 0 640P 0 665P 670U 700P 0 840P 0 865P 670U 900P 0  1040P 0 1065P 670U 1100P 0 1240P 0 1265P 670U 1300P 0  )
LSYNB21 ACTUALSYNB21x ACTUALSYNB21 1p  
KSYNB21 LSYNB21 LSYNADJUSTB21 -0.1
LSYNADJUSTB21 0 ADJUSTB21 5P 

#SPLIT TARGET BETWEEN 2 NEURONS
LTARGET1 TARGET0 TARGET1 1p
LTARGET2 TARGET0 TARGET2 1p

#SPLIT INPUTS BETWEEN 2 NEURONS
LINPUT1 IN1 INPUT11 1P
LINPUT2 IN1 INPUT12 1P
LINPUT3 IN2 INPUT13 1P
LINPUT4 IN2 INPUT14 1P
LINPUTBIAS11 INB11 INPUTB12 1P
LINPUTBIAS12 INB11 INPUTB13 1P


IINITALB21 0 INITIALB21 PWL( 0 0 20P -4*2*22.6U)
XSTOREB21 BISTORE SFQOUTPLUSB21 SFQOUTMINUSB21 WEIGHTLB21 WEIGHTRB21
#IINplusB21 0 INPLUSB21 PULSE(0 000U 2800p 2.5P 2.5P 1P 600P )
#XWEIGHTB21 LSmitll_DCSFQ_PTLTX INPLUSB21 SFQOUTPLUSB21
#IINminusB21 0 INMINUSB21 PULSE(0 000U 400p 2.5P 2.5P 1P 600P )
#IINminusB21cancel21 0 INMINUSB21 PULSE(0 -00U 2200p 2.5P 2.5P 1P 600P )
#XWEIGHTMINUSB21 LSmitll_DCSFQ_PTLTX INMINUSB21 SFQOUTMINUSB21

X21 SYNAPSEfastestnext2 OUTPUTAXON DOUT22 DOUT21  WEIGHTL21 WEIGHTR21 INITIAL21
XB21 SYNAPSEfastestnext2 ACTUALSYNB21  0 DOUT23   WEIGHTLB21 WEIGHTRB21 INITIALB21

IINITAL11 0 INITIAL11 PWL( 0 0 20P -80U)
IINITAL12 0 INITIAL12 PWL( 0 0 20P 0U)
IINITALB11 0 INITIALB11 PWL( 0 0 20P -80U)

IINITAL13 0 INITIAL13 PWL( 0 0 20P -80U)
IINITAL14 0 INITIAL14 PWL( 0 0 20P 0U)
IINITALB12 0 INITIALB12 PWL( 0 0 20P -80U)


##FINAL ACTIVATION - this works 
#ITHRESH11 0 THRESH11 PWL(0 0 20p 200U)
#ITHRESH12 0 THRESH12 PWL(0 0 20p 18U)
#ITHRESH21 0 THRESH21 PWL(0 0 20p -20U)
ITHRESH11 0 THRESH11 PWL(0 0 20p 200U)
ITHRESH12 0 THRESH12 PWL(0 0 20p 200U)
ITHRESH21 0 THRESH21 PWL(0 0 20p 20U)
#was like 23u
XACTfinal COMP6 A5 DOUT21 A6  DC6 DC5   DOUTFINAL1 0   DOUTFINAL2 0   DOUTFINAL3 0  0 DOUTFINAL4   DOUTFINAL5 0 DOUTFINAL6 0   THRESH21

XNEURON1 3NEURON2 INPUT11 INPUT13 INPUTB12 TARGET1 DOUTFINAL1 DOUTFINAL2 THRESH11 A3 A5 B3 B4 DC3 DC5 DCC3 DCC4 OUTPUT1 OUTPUT2 OUTPUTAXON DELAYEDTARGETP DELAYEDTARGETN  DELAYEDTARGETp2 INITIAL11 INITIAL12 INITIALB11
          #x3NEURON2 INPUT1 INPUT2 INPUTBIAS TARGET DOUTFINAL1 DOUTFINAL2 THRESH XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT DCCIN DCCOUT OUTPUT OUTPUTAXON

#xbfrout1 bfr B4 DOUTFINAL3 B5 dc6 DC7  0 actfinaloutp  
xbfrout1 bfrsplit4 B4 DOUTFINAL3 B6 dc6 DC8  0 actfinaloutp  actfinaloutn 0 0 actfinaloutp2  actfinaloutn2 0 
#xbfrout2 bfr B5 DOUTFINAL4 B6 dc7 DC8  0 actfinaloutn 
#xbfrout2 bfrsplit2 B5 DOUTFINAL4 B6 dc7 DC8  0 actfinaloutp2  0 actfinaloutn2 


#xbfrout2 bfr B5 DOUTFINAL4 B6 dc7 DC8  0 actfinaloutn2 actfinaloutp2 0

XPERCEPTRON21 PERCEPTRON   B6  B7 A7 A6   OUTPUT1  actfinaloutp actfinaloutn DELAYEDTARGETP   DC8 DC9 INCR21 DECR21
XCONVO CONV A7 A8   DCC5 DCC4  INCR21 DECR21 SFQOUTPLUS21 SFQOUTMINUS21

XPERCEPTRONb21 PERCEPTRON   B7  B8 A9 A8   ADJUSTB21  actfinaloutp2 actfinaloutn2 DELAYEDTARGETP2   DC9 DC10 INCRb21 DECRb21
XCONVb21 CONV A9 A10   DCC6 DCC5  INCRb21 DECRb21 SFQOUTPLUSb21 SFQOUTMINUSb21

XNEURON2 3NEURON2 INPUT12 INPUT14 INPUTB13 TARGET2 DOUTFINAL5 DOUTFINAL6 THRESH12 A10 A11 B8 B9 DC10 DC11 DCC6 DCC7 OUTPUT3 OUTPUT4 OUTPUTAXON2 DELAYEDTARGETP12 DELAYEDTARGETN12  DELAYEDTARGETP13 INITIAL13 INITIAL14 INITIALB12
IINITAL22 0 INITIAL22 PWL( 0 0 20P -4*2*22.6U)
XSTORE22 BISTORE SFQOUTPLUS22 SFQOUTMINUS22 WEIGHTL22 WEIGHTR22


X22 SYNAPSEfastestnext2 OUTPUTAXON2 DOUT23 DOUT22  WEIGHTL22 WEIGHTR22 INITIAL22
xbfrout2 bfrsplit2 B9 DOUTFINAL4 B10 DC11 DC12 0 actfinaloutp3  actfinaloutn3 0
XPERCEPTRON22 PERCEPTRON   B10  0 A12 A11   OUTPUT3  actfinaloutp3 actfinaloutn3 DELAYEDTARGETP12   DC12 0 INCR22 DECR22
XCONVO22 CONV A12 0   0 DCC7  INCR22 DECR22 SFQOUTPLUS22 SFQOUTMINUS22


#extra set of inputs
#going to need to add another neuron obviously
#another synapse (22)
#buffout3
#perceptron22
#conv22

#XNEURON2 3NEURON2 INPUT13 INPUT14 INB11 TARGET1 DOUTFINAL4 DOUTFINAL5 THRESH11 A3 A5 B3 B4 DC3 DC5 DCC3 DCC4 OUTPUT1 OUTPUT2 OUTPUTAXON DELAYEDTARGETP DELAYEDTARGETN  DELAYEDTARGETp2 INITIAL11 INITIAL12 INITIALB11




.PRINT DEVII IIN1
.PRINT DEVII IIN2
.PRINT DEVII ITARGET
.print devii Iactualsynbias21
.print phase lstore1.x11.XNEURON1
.print phase lstore1.x12.XNEURON1
.print phase lstore1.xb11.XNEURON1
.PRINT PHASE LQ.XACT11.XNEURON1
.PRINT PHASE LQ.XACT11.XNEURON2
.PRINT PHASE LQ.X21
.print phase lstore1.X21
.PRINT PHASE LSTORE1.X22
.print phase lstore1.Xb21
.PRINT PHASE LQ.XACTfinal
.print phase lq.XINPUT.XPERCEPTRON21
.print phase lq.XTARGET.XPERCEPTRON21
.print phase L1_Q.xINCR.XPERCEPTRON21
.print phase L2_Q.xINCR.XPERCEPTRON21
.print phase L4_Q.xINCR.XPERCEPTRON21






.SUBCKT 3NEURON2 INPUT1 INPUT2 INPUTBIAS TARGET ACTNEXT1 ACTNEXT2 THRESH XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT DCCIN DCCOUT OUTPUT1 OUTPUT2 OUTPUTAXON DELAYOUTTARGET3 DELAYOUTTARGET4 DELAYOUTTARGET5 INITIAL11 INITIAL12 INITIALB11

#INPUTS
LSYN11 INPUT1 SYN11 1p  
LSYN12 INPUT2 SYN12 1p  
LSYNB11 INPUTBIAS SYNB11 1p  
LTARGET1 TARGET TARGET1 1p
LTARGET2 TARGET1 0 1p

#COUPLINGS
KSYN11 LSYN11 LSYNADJUST11 -0.05
KSYN12 LSYN12 LSYNADJUST12 -0.05
KSYNB11 LSYNB11 LSYNADJUSTB11 -0.05
KT1 LTARGET1 LADJUSTTARGET1 -0.05
KT2 LTARGET2 LADJUSTTARGET2 -0.05
LSYNADJUST11 0 ADJUST11 5P 
LSYNADJUST12 0 ADJUST12 5P 
LSYNADJUSTB11 0 ADJUSTB11 5P 
LADJUSTTARGET1 0 ADJUSTTARGET1 5P
LADJUSTTARGET2 0 ADJUSTTARGET2 5P


#SYNAPSE 1
#IINITAL11 0 INITIAL11 PWL( 0 0 20P -80U)
XSTORE11 BISTORE SFQOUTPLUS11 SFQOUTMINUS11 WEIGHTL11 WEIGHTR11
X11 SYNAPSEfastest SYN11 DOUT12 DOUT11 WEIGHTL11 WEIGHTR11 INITIAL11
#l111 SFQOUTPLUS11 0 1p
#l112 SFQOUTMINUS11 0 1p

#SYNAPSE 2
#IINITAL12 0 INITIAL12 PWL( 0 0 20P -80U)
XSTORE12 BISTORE SFQOUTPLUS12 SFQOUTMINUS12 WEIGHTL12 WEIGHTR12
X12 SYNAPSEfastest SYN12 DOUT13 DOUT12 WEIGHTL12 WEIGHTR12 INITIAL12
#l121 SFQOUTPLUS12 0 1p
#l122 SFQOUTMINUSB12 0 1p

#SYNAPSE BIAS
#IINITALB11 0 INITIALB11 PWL( 0 0 20P -80U)
XSTOREB11 BISTORE SFQOUTPLUSB11 SFQOUTMINUSB11 WEIGHTLB11 WEIGHTRB11
XB11 SYNAPSEfastest SYNB11 0 DOUT13 WEIGHTLB11 WEIGHTRB11 INITIALB11
#lB111 SFQOUTPLUSB11 0 1p
#lB112 SFQOUTMINUSB11 0 1p

#ACTIVATION
XACT11 COMP5 XIN1 DOUT11 A4 DCIN DC4 DOUTL11 0  0 DOUTR12  0 DOUTL13 0 OUTPUT1 0 OUTPUT2   THRESH

#AXON FOR OUTPUT
XTRANSMIT1 TRANSMIT DOUTL11 XIN2 B4 A4 A6 DC4 DC6 DCCIN DCC4 OUTPUTAXON

#DELAYS
XDELAYACT1 DELAY10 DOUTR12 B4 B5 A6 A7 DC6 DC7  DELAYOUT1 0  DELAYOUT2 0
XDELAYTARGET DELAY14 ADJUSTTARGET1 B5 B6 A7 A8 DC7 DC8   DELAYOUTTARGET1  0 DELAYOUTTARGET2 0


#LEARNING ALGORITHMS
#ASSUME DOUTFINAL1 0 DOUTFINAL2 0  DOUTFINAL3 0  0 DOUTFINAL4
XMLP MLPNEW B6 B7 A8 A9 DELAYOUT1 DELAYOUT2 DELAYOUTTARGET1 DELAYOUTTARGET2 ACTNEXT1 ACTNEXT2 DC8 DC9 OUTPUTTARGET1L 0 OUTPUTTARGET2L 0 OUTPUTTARGET3L 0
XDELAYTARGET2 DELAY18 ADJUSTTARGET2 B7 B8 A9 A10 DC9 dc10  0 DELAYOUTTARGET3  DELAYOUTTARGET4 0  0 DELAYOUTTARGET5 0 
XDELAYINPUT1 DELAY18 ADJUST11  B8  B9  A10 A11 DC10 DC11 DELAYOUTINPUT111 0 DELAYOUTINPUT112 0 DELAYOUTINPUT113 0 DELAYOUTINPUT114 0 DELAYOUTINPUT115 0 DELAYOUTINPUT116 0
XDELAYINPUT2 DELAY18 ADJUST12  B9  B10  A11 A12 DC11 DC12 DELAYOUTINPUT121 0 DELAYOUTINPUT122 0 DELAYOUTINPUT123 0 DELAYOUTINPUT124 0 DELAYOUTINPUT125 0 DELAYOUTINPUT126 0
XDELAYINPUTB1 DELAY18 ADJUSTB11  B10  B11  A12 A13 DC12 DC13 DELAYOUTINPUT1B1 0 DELAYOUTINPUT1B2 0 DELAYOUTINPUT1B3 0 DELAYOUTINPUT1B4 0 DELAYOUTINPUT1B5 0 DELAYOUTINPUT1B6 0

XDELAYact2 DELAY15 DOUTL13  B11 B12  A13 A14 DC13 DC14  DELAYOUTact111 0 0  DELAYOUTact112 DELAYOUTact113 0 0  DELAYOUTact114   DELAYOUTact115  0 0  DELAYOUTact116 


XPERCEPTRON11 PERCEPTRON  B13 B12  A14 A15  DELAYOUTINPUT111 DELAYOUTact111 DELAYOUTact112 OUTPUTTARGET1L DC15 DC14 INCR11 DECR11
XPERCEPTRON12 PERCEPTRON  B14 B13  A15 A16  DELAYOUTINPUT121 DELAYOUTact113 DELAYOUTact114 OUTPUTTARGET2L DC16 DC15 INCR12 DECR12
XPERCEPTRONB11 PERCEPTRON  XOUT2 B14  A16 A17  DELAYOUTINPUT1B1 DELAYOUTact115 DELAYOUTact116 OUTPUTTARGET3L DCOUT DC16 INCRB11 DECRB11

XCONV11 CONV A17 A18 DCC5 DCC4 INCR11 DECR11 SFQOUTPLUS11 SFQOUTMINUS11
XCONV12 CONV A18 A19 DCC6 DCC5 INCR12 DECR12 SFQOUTPLUS12 SFQOUTMINUS12
XCONVB11 CONV A19 XOUT1 DCCOUT DCC6 INCRB11 DECRB11 SFQOUTPLUSB11 SFQOUTMINUSB11

.ENDS 3NEURON2


.SUBCKT MLPNEW XIN1 XOUT1 XIN2 XOUT2 OI1 OI2 T1 T2 OJ1 OJ2 DCIN DCOUT OUTPUTTARGET1L OUTPUTTARGET1R OUTPUTTARGET2L OUTPUTTARGET2R OUTPUTTARGET3L OUTPUTTARGET3R
#Oi.T
Xand1  AND  B7 XIN1  XIN2 A9  OI1 T1 DC9 DCIN  andout1
#Oi.!Oj
Xand2  AND B8 B7 A9 A10 OI2 OJ1 DC10 DC9 andout2
#T.!Oj
Xand3  AND B9 B8 A10 A11 T2 OJ2 DC11 DC10 andout3
#D=Oi.T + Oi.!Oj + T.!Oj 
X3OR OR3 B9 XOUT1 XOUT2 A11   ANDOUT1 ANDOUT2 ANDOUT3 DCOUT DC11  OUTPUTTARGET1L 0 OUTPUTTARGET2L 0 OUTPUTTARGET3L 0
.ENDS MLPNEW













.SUBCKT DELAY10 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 XOUT1  DC15 DC14      DELAYOUT9 0
XDELAY10 bfrsplit2 XOUT2 DELAYOUT9 A10   DC15 DCOUT      OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R
.ends DELAY10

.SUBCKT DELAY11 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR XOUT2 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 bfrsplit2 XOUT1 DELAYOUT10 B9   DCOUT DC16   OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R

.ends DELAY11



.SUBCKT DELAY14 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR A11 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 BFR B10 DELAYOUT10 B9   DC17 DC16   DELAYOUT11 0
XDELAY12 BFR A11 DELAYOUT11 A12   DC17 DC18  DELAYOUT12 0
XDELAY13 BFR B10 DELAYOUT12 XOUT1  DC19 DC18  DELAYOUT13 0
XDELAY14 bfrsplit2 XOUT2 DELAYOUT13 A12  DC19 DCOUT  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R


.ends DELAY14

.SUBCKT DELAY15 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R OUTPUT4L OUTPUT4R OUTPUT5L OUTPUT5R OUTPUT6L OUTPUT6R
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR A11 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 BFR B10 DELAYOUT10 B9   DC17 DC16   DELAYOUT11 0
XDELAY12 BFR A11 DELAYOUT11 A12   DC17 DC18  DELAYOUT12 0
XDELAY13 BFR B10 DELAYOUT12 B11  DC19 DC18  DELAYOUT13 0
XDELAY14 BFR XOUT2 DELAYOUT13 A12  DC19 DC20  DELAYOUT14 0

XDELAY15 bfrsplit6 XOUT1 DELAYOUT14 B11 DCOUT DC20  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R OUTPUT4L OUTPUT4R OUTPUT5L OUTPUT5R OUTPUT6L OUTPUT6R

.ends DELAY15



.SUBCKT DELAY16 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR A11 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 BFR B10 DELAYOUT10 B9   DC17 DC16   DELAYOUT11 0
XDELAY12 BFR A11 DELAYOUT11 A12   DC17 DC18  DELAYOUT12 0
XDELAY13 BFR B10 DELAYOUT12 B11  DC19 DC18  DELAYOUT13 0
XDELAY14 BFR A13 DELAYOUT13 A12  DC19 DC20  DELAYOUT14 0
XDELAY15 BFR XOUT1 DELAYOUT14 B11  DC21 DC20  DELAYOUT15 0
XDELAY16 bfrsplit2 A13 DELAYOUT15 XOUT2  DC21 DCOUT  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R
.ends DELAY16


.SUBCKT DELAY18 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R OUTPUT3L OUTPUT3R
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR A11 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 BFR B10 DELAYOUT10 B9   DC17 DC16   DELAYOUT11 0
XDELAY12 BFR A11 DELAYOUT11 A12   DC17 DC18  DELAYOUT12 0
XDELAY13 BFR B10 DELAYOUT12 B11  DC19 DC18  DELAYOUT13 0
XDELAY14 BFR A13 DELAYOUT13 A12  DC19 DC20  DELAYOUT14 0
XDELAY15 BFR B12 DELAYOUT14 B11  DC21 DC20  DELAYOUT15 0
XDELAY16 BFR A13 DELAYOUT15 A14  DC21 DC22  DELAYOUT16 0
XDELAY17 BFR B12 DELAYOUT16 XOUT1  DC23 DC22  DELAYOUT17 0
XDELAY18 bfrsplit3 XOUT2 DELAYOUT17 A14 DC23 DCOUT  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R  OUTPUT3L OUTPUT3R


.ends DELAY18

***    INPUTS  ***
IIN1 0 IN1 PWL(0 0 20P 0 1.5500e-09 0.0000e+00 1.5550e-09 2.0000e-03 1.6050e-09 2.0000e-03
+ 1.6100e-09 0.0000e+00 3.5500e-09 0.0000e+00 3.5550e-09 2.0000e-03
+ 3.6050e-09 2.0000e-03 3.6100e-09 0.0000e+00 5.5500e-09 0.0000e+00
+ 5.5550e-09 2.0000e-03 5.6050e-09 2.0000e-03 5.6100e-09 0.0000e+00
+ 7.5500e-09 0.0000e+00 7.5550e-09 2.0000e-03 7.6050e-09 2.0000e-03
+ 7.6100e-09 0.0000e+00 9.5500e-09 0.0000e+00 9.5550e-09 2.0000e-03
+ 9.6050e-09 2.0000e-03 9.6100e-09 0.0000e+00 1.1550e-08 0.0000e+00
+ 1.1555e-08 2.0000e-03 1.1605e-08 2.0000e-03 1.1610e-08 0.0000e+00
+ 1.3550e-08 0.0000e+00 1.3555e-08 2.0000e-03 1.3605e-08 2.0000e-03
+ 1.3610e-08 0.0000e+00 1.5550e-08 0.0000e+00 1.5555e-08 2.0000e-03
+ 1.5605e-08 2.0000e-03 1.5610e-08 0.0000e+00 1.7550e-08 0.0000e+00
+ 1.7555e-08 2.0000e-03 1.7605e-08 2.0000e-03 1.7610e-08 0.0000e+00
+ 1.9550e-08 0.0000e+00 1.9555e-08 2.0000e-03 1.9605e-08 2.0000e-03
+ 1.9610e-08 0.0000e+00 2.1550e-08 0.0000e+00 2.1555e-08 2.0000e-03
+ 2.1605e-08 2.0000e-03 2.1610e-08 0.0000e+00 2.3550e-08 0.0000e+00
+ 2.3555e-08 2.0000e-03 2.3605e-08 2.0000e-03 2.3610e-08 0.0000e+00
+ 2.5550e-08 0.0000e+00 2.5555e-08 2.0000e-03 2.5605e-08 2.0000e-03
+ 2.5610e-08 0.0000e+00 2.7550e-08 0.0000e+00 2.7555e-08 2.0000e-03
+ 2.7605e-08 2.0000e-03 2.7610e-08 0.0000e+00 2.9550e-08 0.0000e+00
+ 2.9555e-08 2.0000e-03 2.9605e-08 2.0000e-03 2.9610e-08 0.0000e+00
+ 3.1550e-08 0.0000e+00 3.1555e-08 2.0000e-03 3.1605e-08 2.0000e-03
+ 3.1610e-08 0.0000e+00 3.3550e-08 0.0000e+00 3.3555e-08 2.0000e-03
+ 3.3605e-08 2.0000e-03 3.3610e-08 0.0000e+00 3.5550e-08 0.0000e+00
+ 3.5555e-08 2.0000e-03 3.5605e-08 2.0000e-03 3.5610e-08 0.0000e+00
+ 3.7550e-08 0.0000e+00 3.7555e-08 2.0000e-03 3.7605e-08 2.0000e-03
+ 3.7610e-08 0.0000e+00 3.9550e-08 0.0000e+00 3.9555e-08 2.0000e-03
+ 3.9605e-08 2.0000e-03 3.9610e-08 0.0000e+00 4.1550e-08 0.0000e+00
+ 4.1555e-08 2.0000e-03 4.1605e-08 2.0000e-03 4.1610e-08 0.0000e+00
+ 4.3550e-08 0.0000e+00 4.3555e-08 2.0000e-03 4.3605e-08 2.0000e-03
+ 4.3610e-08 0.0000e+00 4.5550e-08 0.0000e+00 4.5555e-08 2.0000e-03
+ 4.5605e-08 2.0000e-03 4.5610e-08 0.0000e+00 4.7550e-08 0.0000e+00
+ 4.7555e-08 2.0000e-03 4.7605e-08 2.0000e-03 4.7610e-08 0.0000e+00
+ 4.9550e-08 0.0000e+00 4.9555e-08 2.0000e-03 4.9605e-08 2.0000e-03
+ 4.9610e-08 0.0000e+00 5.1550e-08 0.0000e+00 5.1555e-08 2.0000e-03
+ 5.1605e-08 2.0000e-03 5.1610e-08 0.0000e+00 5.3550e-08 0.0000e+00
+ 5.3555e-08 2.0000e-03 5.3605e-08 2.0000e-03 5.3610e-08 0.0000e+00
+ 5.5550e-08 0.0000e+00 5.5555e-08 2.0000e-03 5.5605e-08 2.0000e-03
+ 5.5610e-08 0.0000e+00 5.7550e-08 0.0000e+00 5.7555e-08 2.0000e-03
+ 5.7605e-08 2.0000e-03 5.7610e-08 0.0000e+00 5.9550e-08 0.0000e+00
+ 5.9555e-08 2.0000e-03 5.9605e-08 2.0000e-03 5.9610e-08 0.0000e+00
+ 6.1550e-08 0.0000e+00 6.1555e-08 2.0000e-03 6.1605e-08 2.0000e-03
+ 6.1610e-08 0.0000e+00 6.3550e-08 0.0000e+00 6.3555e-08 2.0000e-03
+ 6.3605e-08 2.0000e-03 6.3610e-08 0.0000e+00 6.5550e-08 0.0000e+00
+ 6.5555e-08 2.0000e-03 6.5605e-08 2.0000e-03 6.5610e-08 0.0000e+00
+ 6.7550e-08 0.0000e+00 6.7555e-08 2.0000e-03 6.7605e-08 2.0000e-03
+ 6.7610e-08 0.0000e+00 6.9550e-08 0.0000e+00 6.9555e-08 2.0000e-03
+ 6.9605e-08 2.0000e-03 6.9610e-08 0.0000e+00 7.1550e-08 0.0000e+00
+ 7.1555e-08 2.0000e-03 7.1605e-08 2.0000e-03 7.1610e-08 0.0000e+00
+ 7.3550e-08 0.0000e+00 7.3555e-08 2.0000e-03 7.3605e-08 2.0000e-03
+ 7.3610e-08 0.0000e+00 7.5550e-08 0.0000e+00 7.5555e-08 2.0000e-03
+ 7.5605e-08 2.0000e-03 7.5610e-08 0.0000e+00 7.7550e-08 0.0000e+00
+ 7.7555e-08 2.0000e-03 7.7605e-08 2.0000e-03 7.7610e-08 0.0000e+00
+ 7.9550e-08 0.0000e+00 7.9555e-08 2.0000e-03 7.9605e-08 2.0000e-03
+ 7.9610e-08 0.0000e+00)
IIN2 0 IN2 PWL(0 0 20P 0 3.5500e-09 0.0000e+00 3.5550e-09 2.0000e-03 3.6050e-09 2.0000e-03
+ 3.6100e-09 0.0000e+00 7.5500e-09 0.0000e+00 7.5550e-09 2.0000e-03
+ 7.6050e-09 2.0000e-03 7.6100e-09 0.0000e+00 1.1550e-08 0.0000e+00
+ 1.1555e-08 2.0000e-03 1.1605e-08 2.0000e-03 1.1610e-08 0.0000e+00
+ 1.5550e-08 0.0000e+00 1.5555e-08 2.0000e-03 1.5605e-08 2.0000e-03
+ 1.5610e-08 0.0000e+00 1.9550e-08 0.0000e+00 1.9555e-08 2.0000e-03
+ 1.9605e-08 2.0000e-03 1.9610e-08 0.0000e+00 2.3550e-08 0.0000e+00
+ 2.3555e-08 2.0000e-03 2.3605e-08 2.0000e-03 2.3610e-08 0.0000e+00
+ 2.7550e-08 0.0000e+00 2.7555e-08 2.0000e-03 2.7605e-08 2.0000e-03
+ 2.7610e-08 0.0000e+00 3.1550e-08 0.0000e+00 3.1555e-08 2.0000e-03
+ 3.1605e-08 2.0000e-03 3.1610e-08 0.0000e+00 3.5550e-08 0.0000e+00
+ 3.5555e-08 2.0000e-03 3.5605e-08 2.0000e-03 3.5610e-08 0.0000e+00
+ 3.9550e-08 0.0000e+00 3.9555e-08 2.0000e-03 3.9605e-08 2.0000e-03
+ 3.9610e-08 0.0000e+00 4.3550e-08 0.0000e+00 4.3555e-08 2.0000e-03
+ 4.3605e-08 2.0000e-03 4.3610e-08 0.0000e+00 4.7550e-08 0.0000e+00
+ 4.7555e-08 2.0000e-03 4.7605e-08 2.0000e-03 4.7610e-08 0.0000e+00
+ 5.1550e-08 0.0000e+00 5.1555e-08 2.0000e-03 5.1605e-08 2.0000e-03
+ 5.1610e-08 0.0000e+00 5.5550e-08 0.0000e+00 5.5555e-08 2.0000e-03
+ 5.5605e-08 2.0000e-03 5.5610e-08 0.0000e+00 5.9550e-08 0.0000e+00
+ 5.9555e-08 2.0000e-03 5.9605e-08 2.0000e-03 5.9610e-08 0.0000e+00
+ 6.3550e-08 0.0000e+00 6.3555e-08 2.0000e-03 6.3605e-08 2.0000e-03
+ 6.3610e-08 0.0000e+00 6.7550e-08 0.0000e+00 6.7555e-08 2.0000e-03
+ 6.7605e-08 2.0000e-03 6.7610e-08 0.0000e+00 7.1550e-08 0.0000e+00
+ 7.1555e-08 2.0000e-03 7.1605e-08 2.0000e-03 7.1610e-08 0.0000e+00
+ 7.5550e-08 0.0000e+00 7.5555e-08 2.0000e-03 7.5605e-08 2.0000e-03
+ 7.5610e-08 0.0000e+00 7.9550e-08 0.0000e+00 7.9555e-08 2.0000e-03
+ 7.9605e-08 2.0000e-03 7.9610e-08 0.0000e+00)
IINBIAS1 0 INB11 pulse(0 0.002 550p 5p 5p 50p 1000p)
ITARGET 0 TARGET0  PWL(0 0 20P 0 3.5500e-09 0.0000e+00 3.5550e-09 2.0000e-03 3.6050e-09 2.0000e-03
+ 3.6100e-09 0.0000e+00 7.5500e-09 0.0000e+00 7.5550e-09 2.0000e-03
+ 7.6050e-09 2.0000e-03 7.6100e-09 0.0000e+00 1.1550e-08 0.0000e+00
+ 1.1555e-08 2.0000e-03 1.1605e-08 2.0000e-03 1.1610e-08 0.0000e+00
+ 1.5550e-08 0.0000e+00 1.5555e-08 2.0000e-03 1.5605e-08 2.0000e-03
+ 1.5610e-08 0.0000e+00 1.9550e-08 0.0000e+00 1.9555e-08 2.0000e-03
+ 1.9605e-08 2.0000e-03 1.9610e-08 0.0000e+00 2.3550e-08 0.0000e+00
+ 2.3555e-08 2.0000e-03 2.3605e-08 2.0000e-03 2.3610e-08 0.0000e+00
+ 2.7550e-08 0.0000e+00 2.7555e-08 2.0000e-03 2.7605e-08 2.0000e-03
+ 2.7610e-08 0.0000e+00 3.1550e-08 0.0000e+00 3.1555e-08 2.0000e-03
+ 3.1605e-08 2.0000e-03 3.1610e-08 0.0000e+00 3.5550e-08 0.0000e+00
+ 3.5555e-08 2.0000e-03 3.5605e-08 2.0000e-03 3.5610e-08 0.0000e+00
+ 3.9550e-08 0.0000e+00 3.9555e-08 2.0000e-03 3.9605e-08 2.0000e-03
+ 3.9610e-08 0.0000e+00 4.3550e-08 0.0000e+00 4.3555e-08 2.0000e-03
+ 4.3605e-08 2.0000e-03 4.3610e-08 0.0000e+00 4.7550e-08 0.0000e+00
+ 4.7555e-08 2.0000e-03 4.7605e-08 2.0000e-03 4.7610e-08 0.0000e+00
+ 5.1550e-08 0.0000e+00 5.1555e-08 2.0000e-03 5.1605e-08 2.0000e-03
+ 5.1610e-08 0.0000e+00 5.5550e-08 0.0000e+00 5.5555e-08 2.0000e-03
+ 5.5605e-08 2.0000e-03 5.5610e-08 0.0000e+00 5.9550e-08 0.0000e+00
+ 5.9555e-08 2.0000e-03 5.9605e-08 2.0000e-03 5.9610e-08 0.0000e+00
+ 6.3550e-08 0.0000e+00 6.3555e-08 2.0000e-03 6.3605e-08 2.0000e-03
+ 6.3610e-08 0.0000e+00 6.7550e-08 0.0000e+00 6.7555e-08 2.0000e-03
+ 6.7605e-08 2.0000e-03 6.7610e-08 0.0000e+00 7.1550e-08 0.0000e+00
+ 7.1555e-08 2.0000e-03 7.1605e-08 2.0000e-03 7.1610e-08 0.0000e+00
+ 7.5550e-08 0.0000e+00 7.5555e-08 2.0000e-03 7.5605e-08 2.0000e-03
+ 7.5610e-08 0.0000e+00 7.9550e-08 0.0000e+00 7.9555e-08 2.0000e-03
+ 7.9605e-08 2.0000e-03 7.9610e-08 0.0000e+00)

#works well!
#got the data to propagate
.include LSmitll_DCSFQ_PTLTX_v1p5.cir
.include LSmitll_PTLRX_SFQDC_v1p5.cir
.include LSmitll_SPLITT_v1p5.cir
.INCLUDE LSMITLL_JTLT_V1P5.CIR
.INCLUDE LSMITLL_MERGET_V1P5.CIR
.include storeedit.cir
.INCLUDE COMPONENTSEDIT.CIR
.INCLUDE COMP3.CIR
.INCLUDE COMP4.CIR
.include conv.cir
.INCLUDE synapsenext2.CIR
.INCLUDE DCPULSER.CIR
.INCLUDE MULTISPLIT.CIR
.include transmit.cir
#.INCLUDE MLP.CIR - USED ONE IN THIS FILE
.INCLUDE DELAY7.CIR
.INCLUDE AND.CIR
.INCLUDE OR3.CIR
.include PERCEPTRON.CIR


# TRY SHIFTING CLK OF OUTPUT BACK A BIT...

.tran 1ps 2000PS 0ps 1p


#setup circuitry
VAC1   A1   0   SIN(0 723mV 10GHz 200Ps 0)
RAC1   A1   A2   1000
LAC1   A2   A3   0.1p
VAC2   B1   0   SIN(0 723mV 10GHz 175.0ps 0)
RAC2   B1   B2   1000
LAC2   B2   B3   0.1p
VDC    DC1   0   pwl(0 0 20p 1023mV)
RDC    DC1   DC2   1000
LDC    DC2   DC3  0.1p
VDCconv    DCc1   0   PWL(0ps 0mV 20ps 1023mV 1.881e-08 1023mV 1.8811000000000002e-08 0)
RDCconv    DCc1   DCc2  640
LDCconv    DCc2   DCc3   0.1p

#need to change inputs now

#############################################INPUTS#####################################################
#Iactualsyn11 0 ACTUALSYN11x PWL(0 0 20P 0 950P 0 955P 1000U)

Iactualsyn11 0 ACTUALSYN11X PWL(0 0 350P 0 550P 0 555P 1000U 605P 1000U 610P 0 750P 0 950P 0 955P 1000U 1005P 1000U 1010P 0 )
Iactualsyn12 0 ACTUALSYN12 PWL(0 0 350P 0 550P 0 555P 0 605P 0 610P 0 750P 0 755P 1000U 805P 1000U 810P 0 950P 0 955P 1000U 1005P 1000U 1010P 0 )
Iactualsynbias11 0 ACTUALSYNB11 PWL(0 0 350P 0 355P 1000U 405P 1000U 410P 0  550P 0 555P 1000U 605P 1000U 610P 0 750P 0 755P 1000U 805P 1000U 810P 0 950P 0 955P 1000U 1005P 1000U 1010P 0 )

#Iactualsyn11 0 ACTUALSYN11 PWL(0 0 395P 0 400P 1000U 450P 1000U 455P 0 600P 0 800P 0 805P 1000U 855P 1000U 860P 0 )
#Iactualsyn12 0 ACTUALSYN12 PWL(0 0 595p 0 600P 1000u 650P 1000U 655P 0 795p 0 800p 1000U 850P 1000u 855P 0 860p 0)
#Iactualsynbias11 0 ACTUALSYNB11 PWL(0 0 250P 0 255P 1000U 305P 1000U 310P 0  450P 0 455P 1000U 505P 1000U 510P 0 650P 0 655P 1000U 705P 1000U 710P 0 850P 0 855P 1000U 905P 1000U 910P 0 )


Iactualsynbias21 0 ACTUALSYNB21 PWL(0 0 640P 0 665P 670U 700P 0 840P 0 865P 670U 900P 0  1040P 0 1065P 670U 1100P 0 1240P 0 1265P 670U 1300P 0  )
#Itarget 0 TARGET0 PWL(0 0 350P 0 550P 0 555P 1000U 605P 1000U 610P 0 750P 0 950P 0 955P 1000U 1005P 1000U 1010P 0 )
ITARGET 0 TARGET0 PWL(0 0 20P 0 950P 0 955P 1000U 1400P 1000U 1401P 0)
LSYN11 ACTUALSYN11X ACTUALSYN11 1p  
LSYN12 ACTUALSYN12X ACTUALSYN12 1p  
LSYNB11 ACTUALSYNB11X ACTUALSYNB11 1p  
#LSYN13 ACTUALSYN13X ACTUALSYN13 1p  
#LSYN14 ACTUALSYN14X ACTUALSYN14 1p  
#LSYNB12 ACTUALSYNB12X ACTUALSYNB12 1p  
LSYNB21 ACTUALSYNB21X ACTUALSYNB21 1p 
LTARGET1 TARGET0 TARGET1 1p
LTARGET2 TARGET1 0 1p

KSYN11 LSYN11 LSYNADJUST11 -0.05
KSYN12 LSYN12 LSYNADJUST12 -0.05
#KSYN13 LSYN13 LSYNADJUST13 -0.05
#KSYN14 LSYN14 LSYNADJUST14 -0.05
KSYNB11 LSYNB11 LSYNADJUSTB11 -0.05
#KSYNB12 LSYNB12 LSYNADJUSTB12 -0.05
KSYNB21 LSYNB21 LSYNADJUSTB21 -0.05
KT1 LTARGET1 LADJUSTTARGET1 -0.05
KT2 LTARGET2 LADJUSTTARGET2 -0.05

LSYNADJUST11 0 ADJUST11 5P 
LSYNADJUST12 0 ADJUST12 5P 
#LSYNADJUST13 0 ADJUST13 5P 
#LSYNADJUST14 0 ADJUST14 5P 
LSYNADJUSTB11 0 ADJUSTB11 5P 
#LSYNADJUSTB12 0 ADJUSTB12 5P 
LSYNADJUSTB21 0 ADJUSTB21 5P 
LADJUSTTARGET1 0 ADJUSTTARGET1 5P
LADJUSTTARGET2 0 ADJUSTTARGET2 5P

##################################################################

#NEURON1#####################

#SYNAPSE 1 SETUP
#Iactualsyn11 0 ACTUALSYN11 PWL(0 0 350P 0 550P 0 555P 1000U 605P 1000U 610P 0 750P 0 950P 0 955P 1000U 1005P 1000U 1010P 0 )
IINITAL11 0 INITIAL11 PWL( 0 0 20P -80U)
XSTORE11 BISTORE SFQOUTPLUS11 SFQOUTMINUS11 WEIGHTL11 WEIGHTR11
IINplus11 0 INPLUS11 PULSE(0 00U 2800p 2.5P 2.5P 1P 600P )
#IINplus1cancel 0 INPLUS11 PULSE(0 00U 400p 2.5P 2.5P 1P 600P )
XWEIGHT11 LSmitll_DCSFQ_PTLTX INPLUS11 SFQOUTPLUS11
IINminus11 0 INMINUS11 PULSE(0 00U 400p 2.5P 2.5P 1P 600P )
IINminus1cancel11 0 INMINUS11 PULSE(0 -00U 2200p 2.5P 2.5P 1P 600P )
XWEIGHTMINUS11 LSmitll_DCSFQ_PTLTX INMINUS11 SFQOUTMINUS11

#SYNAPSE 2 setup
#Iactualsyn12 0 ACTUALSYN12 PWL(0 0 350P 0 550P 0 555P 0 605P 0 610P 0 750P 0 755P 1000U 805P 1000U 810P 0 950P 0 955P 1000U 1005P 1000U 1010P 0 )

IINITAL12 0 INITIAL12 PWL( 0 0 20P -80U)
XSTORE12 BISTORE SFQOUTPLUS12 SFQOUTMINUS12 WEIGHTL12 WEIGHTR12
IINplus12 0 INPLUS12 PULSE(0 00U 2800p 2.5P 2.5P 1P 600P )
XWEIGHT12 LSmitll_DCSFQ_PTLTX INPLUS12 SFQOUTPLUS12
IINminus12 0 INMINUS12 PULSE(0 00U 400p 2.5P 2.5P 1P 600P )
IINminus2cancel12 0 INMINUS12 PULSE(0 -000U 2200p 2.5P 2.5P 1P 600P )
XWEIGHTMINUS12 LSmitll_DCSFQ_PTLTX INMINUS12 SFQOUTMINUS12


#SYNAPSE bias 1 setup
#IactualsynBIAS11 0 ACTUALSYNB11 PWL(0 0 350P 0 355P 1000U 405P 1000U 410P 0  550P 0 555P 1000U 605P 1000U 610P 0 750P 0 755P 1000U 805P 1000U 810P 0 950P 0 955P 1000U 1005P 1000U 1010P 0 )

IINITALB11 0 INITIALB11 PWL( 0 0 20P -80U)
XSTOREB11 BISTORE SFQOUTPLUSB11 SFQOUTMINUSB11 WEIGHTLB11 WEIGHTRB11
IINplusB11 0 INPLUSB11 PULSE(0 000U 2800p 2.5P 2.5P 1P 600P )
XWEIGHTB11 LSmitll_DCSFQ_PTLTX INPLUSB11 SFQOUTPLUSB11
IINminusB11 0 INMINUSB11 PULSE(0 000U 400p 2.5P 2.5P 1P 600P )
IINminusBcancel11 0 INMINUSB11 PULSE(0 -000U 2200p 2.5P 2.5P 1P 600P )
XWEIGHTMINUSB11 LSmitll_DCSFQ_PTLTX INMINUSB11 SFQOUTMINUSB11

#SYNAPSES FIRST LAYER 1
X11 SYNAPSEfastest ACTUALSYN11 DOUT12 DOUT11 WEIGHTL11 WEIGHTR11 INITIAL11
X12 SYNAPSEfastest ACTUALSYN12 DOUT13 DOUT12 WEIGHTL12 WEIGHTR12 INITIAL12
XB11 SYNAPSEfastest ACTUALSYNB11 0 DOUT13 WEIGHTLB11 WEIGHTRB11 INITIALB11

#ACTIVATION
ITHRESH11 0 THRESH11 PWL(0 0 20p 34U)
#WAS 22
#25 worsk

#TRIED DOUBLING CLK
#XACT11 COMP3 A3 DOUT11 A4 DC3 DC4 DOUTL11 0  DOUTL12 0 0 DOUTL13 THRESH11
XACT11 COMP4 A3 DOUT11 A4 DC3 DC4 DOUTL11 0  0 DOUTR12  0 DOUTL13 DOUTL14 0  THRESH11


##NEURON2#####################



#TRANSMISISON STAGE
XTRANSMIT1 TRANSMIT DOUTL11 B3 B4 A4 A5 DC4 DC5 DCc3 0 OUTCOMBINED11

#XTRANSMIT1 TRANSMIT DOUTL11 B3 0 A5 A6 DC5 DC6 DCc3 DCc4 OUTCOMBINED11
#XTRANSMIT2 TRANSMIT DOUTL14 B4 0 A6 A7 DC6 DC7 DCc4 0 OUTCOMBINED12


#SECOND LAYER SYNAPSE 1

IINITAL21 0 INITIAL21 PWL( 0 0 20P 3*2*22.6U)
XSTORE21 BISTORE SFQOUTPLUS21 SFQOUTMINUS21 WEIGHTL21 WEIGHTR21
IINplusN21 0 INPLUS21 PULSE(0 00U 7400p 2.5P 2.5P 1P 600P )
IINPLUS21cancel21 0 INPLUS21 PULSE(0 -600U 11000p 2.5P 2.5P 1P 600P )
XWEIGHT21 LSmitll_DCSFQ_PTLTX INPLUS21 SFQOUTPLUS21
IINminus21 0 INMINUS21 PULSE(0 00U 11000p 2.5P 2.5P 1P 600P )
IINminuscancel21 0 INMINUS21 PULSE(0 -00U 2800p 2.5P 2.5P 1P 600P )
XWEIGHTMINUS21 LSmitll_DCSFQ_PTLTX INMINUS21 SFQOUTMINUS21

#NEXT LAYER BIAS
#Iactualsynbias21 0 ACTUALSYNB21 PWL(0 0 640P 0 665P 670U 700P 0 840P 0 865P 670U 900P 0  1040P 0 1065P 670U 1100P 0 1240P 0 1265P 670U 1300P 0  )
IINITALB21 0 INITIALB21 PWL( 0 0 20P -4*2*22.6U)
XSTOREB21 BISTORE SFQOUTPLUSB21 SFQOUTMINUSB21 WEIGHTLB21 WEIGHTRB21
IINplusB21 0 INPLUSB21 PULSE(0 000U 2800p 2.5P 2.5P 1P 600P )
XWEIGHTB21 LSmitll_DCSFQ_PTLTX INPLUSB21 SFQOUTPLUSB21
IINminusB21 0 INMINUSB21 PULSE(0 000U 400p 2.5P 2.5P 1P 600P )
IINminusB21cancel21 0 INMINUSB21 PULSE(0 -00U 2200p 2.5P 2.5P 1P 600P )
XWEIGHTMINUSB21 LSmitll_DCSFQ_PTLTX INMINUSB21 SFQOUTMINUSB21


#SECOND LAYER SYNAPSES
#SWITCHED OUTPUT POLARITY
X21 SYNAPSEfastestnext2 OUTCOMBINED11 DOUT23 DOUT21  WEIGHTL21 WEIGHTR21 INITIAL21
#X22 SYNAPSEfastestnext2 OUTCOMBINED12 DOUT23 DOUT22  WEIGHTL22 WEIGHTR22 INITIAL22
XB21 SYNAPSEfastestnext2 ACTUALSYNB21  0 DOUT23   WEIGHTLB21 WEIGHTRB21 INITIALB21

##FINAL ACTIVATION - this works 

#ITHRESH21 0 THRESH21 PWL(0 0 20p -20U)
#XACTfinal COMP3 0 DOUT21 C3  0 DC7  DOUTfinal1 0  DOUTfinal2 0 0 DOUTfinal3 THRESH21
ITHRESH21 0 THRESH21 PWL(0 0 20p -20U)
#was like 23u
XACTfinal COMP3 A5 DOUT21 A6  DC6 DC5  DOUTFINAL1 0   DOUTFINAL2 0  DOUTFINAL3 0 THRESH21

#ACTIVATION, TARGET OUTPUT
#XMLP MLP DOUTR2 ADJUSTTARGET DOUTFINAL1 DOUTLFINAL2 B4 0 A6 0 DC6 0 0 OUTPUTTARGET1R 0 OUTPUTTARGET2R

XDELAYACT1 DELAY10 DOUTR12 B4 B5 A6 A7 DC6 DC7  DELAYOUT1 0  DELAYOUT2 0
XDELAYTARGET DELAY14 ADJUSTTARGET1 B5 B6 A7 A8 DC7 DC8   DELAYOUTTARGET1  0 DELAYOUTTARGET2 0



#Xand1  AND  B7 B6  A8 A9  DELAYOUT1 DELAYOUTTARGET1 DC9 DC8  andout1
#Xand2  AND B8 B7 A9 A10 DELAYOUT2 DOUTFINAL1 DC10 DC9 andout2
#Xand3  AND B9 B8 A10 A11 DELAYOUTTARGET2 DOUTFINAL2 DC11 DC10 andout3
##Oi.T + Oi.!Oj + T.!Oj - 
#X3OR OR3 B9 0 0 A11   ANDOUT1 ANDOUT2 ANDOUT3 0 DC11  OUTPUTTARGET1L 0 OUTPUTTARGET2L 0

XMLP MLPNEW B6 B7 A8 A9 DELAYOUT1 DELAYOUT2 DELAYOUTTARGET1 DELAYOUTTARGET2 DOUTFINAL1 DOUTFINAL2 DC8 DC9 OUTPUTTARGET1L 0 OUTPUTTARGET2L 0
#NOW DELAY STUFF SO THAT THEY CAN WORK WITH THE MLP FOR ADJUSTMENT OF SYNAPSE
#DELAY BY A LITTLE MORE
XDELAYTARGET2 DELAY18 ADJUSTTARGET2 B7 B8 A9 A10 DC9 dc10  DELAYOUTTARGET3 0 DELAYOUTTARGET4 0
XDELAYINPUT DELAY18 ADJUST11  B8  B9  A10 A11 DC10 DC11 DELAYOUTINPUT111 0 DELAYOUTINPUT112 0
XDELAYact2 DELAY15 DOUTL13  B9 B10  A11 A12 DC11 DC12 DELAYOUTact111 0 0 DELAYOUTact112 


#check that it works with perceptron ALGORITHM:
#XPERCEPTRON11 AND3  0 B9 A11 0 DELAYOUTTARGET3 delayout



#now first apply PERCEPTRON to output layer:
#!Tox and T!ox
#XINCR21 AND3  0 B9 A11 0 DELAYOUTTARGET3 doutfinal3 
#XPERCEPTRON11 PERCEPTRON 0 B10 A12 0 DELAYOUTINPUT111 DELAYOUTact111 DELAYOUTact112 OUTPUTTARGET1L 0 DC12 INCR DECR
XPERCEPTRON11 PERCEPTRON  0 B10  A12 0  DELAYOUTINPUT111 DELAYOUTact111 DELAYOUTact112 OUTPUTTARGET1L 0 DC12 INCR DECR



LT1 ADJUST11 0 5p
.print devii Iactualsyn11
.print devii Iactualsyn12
.PRINT DEVII Itarget
.print devii Iactualsynbias11
.print PHASE lq.XACT11
.print devii lstore1.X21
#.print phase b1.X21
#.print phase b2.x21
#.print nodep left.x21
#.print nodep right.x21
.PRINT PHASE LQ.X21
#.PRINT phase LQ.XB21
.PRINT PHASE LQ.XACTfinal
#.print PHASE LQ.XDELAY10.XDELAYACT1
#.print PHASE LQ.XDELAY14.XDELAYTARGET
#.PRINT PHASE L4_Q.XAND1.XMLP
#.PRINT PHASE L4_Q.XAND2.XMLP
#.PRINT PHASE L4_Q.XAND3.XMLP
#.PRINT PHASE L1_Q.X3OR.XMLP
#.PRINT PHASE L2_Q.X3OR.XMLP
#.PRINT PHASE L4_Q.X3OR.XMLP
.PRINT PHASE L5_Q.X3OR.XMLP
.print phase lq.XDELAY15.XDELAYACT2
.PRINT PHASE LQ.XINPUT.XPERCEPTRON11
#.PRINT PHASE LQ.XTARGET.XPERCEPTRON11
.PRINT PHASE L5_Q.XINCR.XPERCEPTRON11
.PRINT PHASE L5_Q.XDECR.XPERCEPTRON11

#.PRINT PHASE L1_Q.XINCR.XPERCEPTRON11
#.PRINT PHASE L2_Q.XINCR.XPERCEPTRON11
#.PRINT PHASE L3_Q.XINCR.XPERCEPTRON11
#.PRINT PHASE L4_Q.XINCR.XPERCEPTRON11
#.PRINT PHASE L5_Q.XINCR.XPERCEPTRON11














.SUBCKT DELAY10 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 XOUT1  DC15 DC14      DELAYOUT9 0
XDELAY10 bfrsplit2 XOUT2 DELAYOUT9 A10   DC15 DCOUT      OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R
.ends DELAY10

.SUBCKT DELAY11 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR XOUT2 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 bfrsplit2 XOUT1 DELAYOUT10 B9   DCOUT DC16   OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R

.ends DELAY11



.SUBCKT DELAY14 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR A11 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 BFR B10 DELAYOUT10 B9   DC17 DC16   DELAYOUT11 0
XDELAY12 BFR A11 DELAYOUT11 A12   DC17 DC18  DELAYOUT12 0
XDELAY13 BFR B10 DELAYOUT12 XOUT1  DC19 DC18  DELAYOUT13 0
XDELAY14 bfrsplit2 XOUT2 DELAYOUT13 A12  DC19 DCOUT  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R


.ends DELAY14

.SUBCKT DELAY15 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR A11 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 BFR B10 DELAYOUT10 B9   DC17 DC16   DELAYOUT11 0
XDELAY12 BFR A11 DELAYOUT11 A12   DC17 DC18  DELAYOUT12 0
XDELAY13 BFR B10 DELAYOUT12 B11  DC19 DC18  DELAYOUT13 0
XDELAY14 BFR XOUT2 DELAYOUT13 A12  DC19 DC20  DELAYOUT14 0

XDELAY15 bfrsplit2 XOUT1 DELAYOUT14 B11 DCOUT DC20  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R


.ends DELAY15



.SUBCKT DELAY16 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR A11 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 BFR B10 DELAYOUT10 B9   DC17 DC16   DELAYOUT11 0
XDELAY12 BFR A11 DELAYOUT11 A12   DC17 DC18  DELAYOUT12 0
XDELAY13 BFR B10 DELAYOUT12 B11  DC19 DC18  DELAYOUT13 0
XDELAY14 BFR A13 DELAYOUT13 A12  DC19 DC20  DELAYOUT14 0
XDELAY15 BFR XOUT1 DELAYOUT14 B11  DC21 DC20  DELAYOUT15 0
XDELAY16 bfrsplit2 A13 DELAYOUT15 XOUT2  DC21 DCOUT  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R
.ends DELAY16


.SUBCKT DELAY18 INPUT XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R
XDELAY1 BFR XIN1 INPUT B5 DC7  DCIN  DELAYOUT1 0
XDELAY2 BFR A7 DELAYOUT1 XIN2 DC7 DC8   DELAYOUT2 0
XDELAY3 BFR B6 DELAYOUT2 B5 DC9 DC8   DELAYOUT3 0
XDELAY4 BFR A7 DELAYOUT3 A8 DC9 dc10    DELAYOUT4 0
XDELAY5 BFR B6 DELAYOUT4 B7 DC11 DC10    DELAYOUT5 0
XDELAY6 BFR A9 DELAYOUT5 A8 DC11 DC12    DELAYOUT6 0
XDELAY7 BFR B8 DELAYOUT6 B7  DC13 DC12     DELAYOUT7 0
XDELAY8 BFR A9 DELAYOUT7 A10  DC13 DC14     DELAYOUT8 0
XDELAY9 BFR B8 DELAYOUT8 B9  DC15 DC14      DELAYOUT9 0
XDELAY10 BFR A11 DELAYOUT9 A10   DC15 DC16   DELAYOUT10 0
XDELAY11 BFR B10 DELAYOUT10 B9   DC17 DC16   DELAYOUT11 0
XDELAY12 BFR A11 DELAYOUT11 A12   DC17 DC18  DELAYOUT12 0
XDELAY13 BFR B10 DELAYOUT12 B11  DC19 DC18  DELAYOUT13 0
XDELAY14 BFR A13 DELAYOUT13 A12  DC19 DC20  DELAYOUT14 0
XDELAY15 BFR B12 DELAYOUT14 B11  DC21 DC20  DELAYOUT15 0
XDELAY16 BFR A13 DELAYOUT15 A14  DC21 DC22  DELAYOUT16 0
XDELAY17 BFR B12 DELAYOUT16 XOUT1  DC23 DC22  DELAYOUT17 0
XDELAY18 bfrsplit2 XOUT2 DELAYOUT17 A14 DC23 DCOUT  OUTPUT1L OUTPUT1R OUTPUT2L OUTPUT2R


.ends DELAY18

.subckt MLP ACTIVATIONPREV1 ACTIVATIONPREV2 TARGET1 TARGET2 ACTIVATIONNEXT1 ACTIVATIONNEXT2 XIN1 XOUT1 XIN2 XOUT2 DCIN DCOUT OUTPUTTARGET1L OUTPUTTARGET1R OUTPUTTARGET2L OUTPUTTARGET2R

#need Oi.T + Oi.!Oj + T.!Oj
#delays so timing matches up
#Xactdelayed DELAY7 ACTIVATIONPREV  XIN1 B6 XIN2 A5 DCIN DC6  0 DELAYOUTACT1  0 DELAYOUTACT2
#XTARGETdelayed DELAY7 TARGET  B6 B7 A5 A6 DC6 DC7 0 DELAYOUTTARGET1  0 DELAYOUTTARGET2 

#Oi.T - correct
Xand1  AND XIN1 A7 XIN2 B8 TARGET1 ACTIVATIONPREV1 DCIN DC8 andout1
#Oi.Oj! - correct
Xand2  AND A7 A8 B8 B9 ACTIVATIONPREV2 ACTIVATIONNEXT1 DC8 DC9 andout2
#T.Oj - correct
Xand3  AND A8 A9 B9 B10 TARGET2 ACTIVATIONNEXT2 DC9 DC10 andout3

#MLP : D = Oi.T + Oi.!Oj + T.!Oj - correct
X3OR OR3 XOUT2 A9 XOUT1 B10  ANDOUT1 ANDOUT2 ANDOUT3 DC10 DCOUT OUTPUTTARGET1L OUTPUTTARGET1R OUTPUTTARGET2L OUTPUTTARGET2R

.ends MLP



.SUBCKT MLPNEW XIN1 XOUT1 XIN2 XOUT2 OI1 OI2 T1 T2 OJ1 OJ2 DCIN DCOUT OUTPUTTARGET1L OUTPUTTARGET1R OUTPUTTARGET2L OUTPUTTARGET2R
#Oi.T
Xand1  AND  B7 XIN1  XIN2 A9  OI1 T1 DC9 DCIN  andout1
#Oi.!Oj
Xand2  AND B8 B7 A9 A10 OI2 OJ1 DC10 DC9 andout2
#T.!Oj
Xand3  AND B9 B8 A10 A11 T2 OJ2 DC11 DC10 andout3
#D=Oi.T + Oi.!Oj + T.!Oj 
X3OR OR3 B9 XOUT1 XOUT2 A11   ANDOUT1 ANDOUT2 ANDOUT3 DCOUT DC11  OUTPUTTARGET1L 0 OUTPUTTARGET2L 0
.ENDS MLPNEW

#2.91E-16Wb=-0.88rad
#@1.264ns
#j1 = -2.26
#j2 = 1.2
#phasesum=0.53
#phasedoff=-1.73
#phix-phasesum=0.35
#measure = -0.5

#using nodep:
#2.91E-16Wb=-0.88rad
#@1.264ns
#j1 node = -2.28
#j2 = 1.3
#phasesum=0.49
#phasedoff=-1.79
#phix-phasesum=0.35
#measure = -0.5

#looks like phase across LQ is simply equal to phase sum of the junctions (use nodes to take parasitics into account)